magic
tech scmos
timestamp 1485907293
use inv_4x  inv_4x_0
timestamp 1485568577
transform 1 0 0 0 1 4
box -6 -4 18 96
use nand2_2x  nand2_2x_0
timestamp 1485568973
transform 1 0 30 0 1 4
box -6 -4 26 96
use nor2_2x  nor2_2x_0
timestamp 1485568973
transform 1 0 68 0 1 4
box -6 -4 26 96
use nand3_1_5x  nand3_1_5x_0
timestamp 1485569183
transform 1 0 106 0 1 4
box -6 -4 34 96
use a2o1i_1_5x  a2o1i_1_5x_0
timestamp 1485569429
transform 1 0 150 0 1 4
box -4 -4 36 96
use flop_dp_4x  flop_dp_4x_0
timestamp 1485645272
transform 1 0 158 0 1 4
box 34 -4 146 96
use mux2i_dp_1_5x  mux2i_dp_1_5x_0
timestamp 1485569944
transform 1 0 316 0 1 4
box -6 -4 42 96
<< end >>
