magic
tech scmos
timestamp 1491509845
<< nwell >>
rect -6 40 58 96
<< ntransistor >>
rect 8 8 10 14
rect 16 8 18 22
rect 21 8 23 22
rect 29 8 31 22
rect 34 8 36 22
rect 42 8 44 14
<< ptransistor >>
rect 8 73 10 82
rect 16 62 18 82
rect 21 62 23 82
rect 29 62 31 82
rect 34 62 36 82
rect 42 73 44 82
<< ndiffusion >>
rect 3 13 8 14
rect 7 9 8 13
rect 3 8 8 9
rect 10 8 11 14
rect 15 8 16 22
rect 18 8 21 22
rect 23 17 29 22
rect 23 8 24 17
rect 28 8 29 17
rect 31 8 34 22
rect 36 8 37 22
rect 41 8 42 14
rect 44 13 49 14
rect 44 9 45 13
rect 44 8 49 9
<< pdiffusion >>
rect 7 73 8 82
rect 10 73 11 82
rect 15 62 16 82
rect 18 62 21 82
rect 23 62 24 82
rect 28 62 29 82
rect 31 62 34 82
rect 36 62 37 82
rect 41 73 42 82
rect 44 73 45 82
<< ndcontact >>
rect 3 9 7 13
rect 11 8 15 22
rect 24 8 28 17
rect 37 8 41 22
rect 45 9 49 13
<< pdcontact >>
rect 3 73 7 82
rect 11 62 15 82
rect 24 62 28 82
rect 37 62 41 82
rect 45 73 49 82
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
rect 40 -2 44 2
rect 48 -2 52 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
rect 32 88 36 92
rect 40 88 44 92
rect 48 88 52 92
<< polysilicon >>
rect 8 82 10 84
rect 16 82 18 84
rect 21 82 23 84
rect 29 82 31 84
rect 34 82 36 84
rect 42 82 44 84
rect 8 72 10 73
rect 2 70 10 72
rect 2 42 4 70
rect 42 72 44 73
rect 42 70 49 72
rect 16 61 18 62
rect 10 59 18 61
rect 10 58 12 59
rect 2 17 4 38
rect 9 25 11 38
rect 9 23 18 25
rect 16 22 18 23
rect 21 22 23 62
rect 29 50 31 62
rect 34 57 36 62
rect 47 58 49 70
rect 34 55 42 57
rect 29 22 31 46
rect 40 42 42 55
rect 40 25 42 29
rect 34 23 42 25
rect 34 22 36 23
rect 2 15 10 17
rect 8 14 10 15
rect 47 17 49 54
rect 42 15 49 17
rect 42 14 44 15
rect 8 6 10 8
rect 16 6 18 8
rect 21 6 23 8
rect 29 6 31 8
rect 34 6 36 8
rect 42 6 44 8
<< polycontact >>
rect 8 54 12 58
rect 17 51 21 55
rect 0 38 4 42
rect 8 38 12 42
rect 28 46 32 50
rect 46 54 50 58
rect 39 38 43 42
rect 39 29 43 33
<< metal1 >>
rect -2 92 54 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 32 92
rect 36 88 40 92
rect 44 88 48 92
rect 52 88 54 92
rect -2 86 54 88
rect 11 82 15 86
rect 37 82 41 86
rect 4 54 8 58
rect 17 55 40 58
rect 21 54 40 55
rect 44 54 46 58
rect 32 46 48 50
rect 4 38 8 42
rect 12 38 39 42
rect 4 29 39 33
rect 4 13 7 14
rect 3 8 7 9
rect 24 17 28 22
rect 45 13 48 14
rect 45 8 49 9
rect 11 4 15 8
rect 37 4 41 8
rect -2 2 54 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 40 2
rect 44 -2 48 2
rect 52 -2 54 2
rect -2 -4 54 -2
<< m2contact >>
rect 0 73 3 77
rect 3 73 4 77
rect 24 62 28 66
rect 48 73 49 77
rect 49 73 52 77
rect 0 54 4 58
rect 40 54 44 58
rect 48 46 52 50
rect 8 38 12 42
rect 0 29 4 33
rect 0 13 4 14
rect 0 10 3 13
rect 3 10 4 13
rect 48 13 52 14
rect 48 10 49 13
rect 49 10 52 13
<< metal2 >>
rect 0 58 4 73
rect 0 42 4 54
rect 0 38 3 42
rect 0 33 4 38
rect 0 14 4 29
rect 24 18 28 62
rect 48 50 52 73
rect 48 14 52 46
<< labels >>
rlabel m2contact 10 40 10 40 1 a
rlabel m2contact 42 56 42 56 1 b
rlabel m2contact 26 64 26 64 1 y
<< end >>
