magic
tech scmos
timestamp 1485645272
<< nwell >>
rect 34 40 146 96
<< ntransistor >>
rect 45 8 47 14
rect 61 8 63 14
rect 69 8 71 12
rect 76 8 78 12
rect 85 8 87 14
rect 93 8 95 14
rect 101 8 103 12
rect 108 8 110 12
rect 117 8 119 14
rect 133 7 135 34
<< ptransistor >>
rect 45 71 47 83
rect 61 77 63 83
rect 69 79 71 83
rect 76 79 78 83
rect 85 74 87 83
rect 93 77 95 83
rect 101 79 103 83
rect 108 79 110 83
rect 117 74 119 83
rect 133 46 135 83
<< ndiffusion >>
rect 44 8 45 14
rect 47 8 48 14
rect 60 8 61 14
rect 63 8 64 14
rect 80 13 85 14
rect 68 8 69 12
rect 71 8 76 12
rect 78 9 80 12
rect 84 9 85 13
rect 78 8 85 9
rect 87 8 88 14
rect 92 8 93 14
rect 95 8 96 14
rect 128 32 133 34
rect 100 8 101 12
rect 103 8 108 12
rect 110 8 112 12
rect 116 8 117 14
rect 119 8 120 14
rect 132 8 133 32
rect 128 7 133 8
rect 135 32 140 34
rect 135 8 136 32
rect 135 7 140 8
<< pdiffusion >>
rect 44 71 45 83
rect 47 71 48 83
rect 60 77 61 83
rect 63 77 64 83
rect 68 79 69 83
rect 71 79 76 83
rect 78 79 80 83
rect 84 74 85 83
rect 87 74 88 83
rect 92 77 93 83
rect 95 77 96 83
rect 100 79 101 83
rect 103 79 108 83
rect 110 79 112 83
rect 116 74 117 83
rect 119 74 120 83
rect 128 81 133 83
rect 132 47 133 81
rect 128 46 133 47
rect 135 81 140 83
rect 135 47 136 81
rect 135 46 140 47
<< ndcontact >>
rect 40 8 44 14
rect 48 8 52 14
rect 56 8 60 14
rect 64 8 68 14
rect 80 9 84 13
rect 88 8 92 14
rect 96 8 100 14
rect 112 8 116 14
rect 120 8 124 14
rect 128 8 132 32
rect 136 8 140 32
<< pdcontact >>
rect 40 71 44 83
rect 48 71 52 83
rect 56 77 60 83
rect 64 77 68 83
rect 80 74 84 83
rect 88 74 92 83
rect 96 77 100 83
rect 112 74 116 83
rect 120 74 124 83
rect 128 47 132 81
rect 136 47 140 81
<< psubstratepcontact >>
rect 40 -2 44 2
rect 48 -2 52 2
rect 56 -2 60 2
rect 64 -2 68 2
rect 72 -2 76 2
rect 80 -2 84 2
rect 88 -2 92 2
rect 96 -2 100 2
rect 104 -2 108 2
rect 112 -2 116 2
rect 120 -2 124 2
rect 128 -2 132 2
rect 136 -2 140 2
<< nsubstratencontact >>
rect 40 88 44 92
rect 48 88 52 92
rect 56 88 60 92
rect 64 88 68 92
rect 72 88 76 92
rect 80 88 84 92
rect 88 88 92 92
rect 96 88 100 92
rect 104 88 108 92
rect 112 88 116 92
rect 120 88 124 92
rect 128 88 132 92
rect 136 88 140 92
<< polysilicon >>
rect 45 83 47 85
rect 61 83 63 85
rect 69 83 71 85
rect 76 83 78 85
rect 85 83 87 85
rect 93 83 95 85
rect 101 83 103 85
rect 108 83 110 85
rect 117 83 119 85
rect 133 83 135 85
rect 45 47 47 71
rect 61 57 63 77
rect 69 74 71 79
rect 76 67 78 79
rect 76 63 77 67
rect 61 45 63 53
rect 61 43 71 45
rect 45 14 47 43
rect 61 14 63 17
rect 69 12 71 43
rect 76 12 78 63
rect 85 28 87 74
rect 93 57 95 77
rect 101 74 103 79
rect 108 67 110 79
rect 108 63 109 67
rect 96 53 103 55
rect 86 24 87 28
rect 85 14 87 24
rect 93 14 95 17
rect 101 12 103 53
rect 108 12 110 63
rect 117 36 119 74
rect 118 32 119 36
rect 133 34 135 46
rect 117 14 119 32
rect 45 6 47 8
rect 61 6 63 8
rect 69 6 71 8
rect 76 6 78 8
rect 85 6 87 8
rect 93 6 95 8
rect 101 6 103 8
rect 108 6 110 8
rect 117 6 119 8
rect 133 5 135 7
<< polycontact >>
rect 68 70 72 74
rect 77 63 81 67
rect 60 53 64 57
rect 44 43 48 47
rect 60 17 64 21
rect 100 70 104 74
rect 109 63 113 67
rect 92 53 96 57
rect 82 24 86 28
rect 92 17 96 21
rect 129 39 133 43
rect 114 32 118 36
<< metal1 >>
rect 38 92 142 94
rect 38 88 40 92
rect 44 88 48 92
rect 52 88 56 92
rect 60 88 64 92
rect 68 88 72 92
rect 76 88 80 92
rect 84 88 88 92
rect 92 88 96 92
rect 100 88 104 92
rect 108 88 112 92
rect 116 88 120 92
rect 124 88 128 92
rect 132 88 136 92
rect 140 88 142 92
rect 38 86 142 88
rect 40 83 44 86
rect 80 83 84 86
rect 112 83 116 86
rect 56 74 60 77
rect 52 71 56 74
rect 48 70 56 71
rect 88 67 92 74
rect 120 67 124 74
rect 81 63 88 67
rect 113 63 124 67
rect 64 53 80 57
rect 96 53 112 57
rect 120 43 124 63
rect 128 81 132 86
rect 128 46 132 47
rect 136 81 140 83
rect 136 46 140 47
rect 124 39 129 43
rect 48 30 56 34
rect 100 32 114 36
rect 128 32 132 34
rect 48 14 52 30
rect 68 24 82 28
rect 104 21 108 25
rect 64 17 72 21
rect 96 17 108 21
rect 80 13 84 14
rect 40 4 44 8
rect 80 4 84 9
rect 112 4 116 8
rect 128 4 132 8
rect 136 32 140 42
rect 136 7 140 8
rect 38 2 142 4
rect 38 -2 40 2
rect 44 -2 48 2
rect 52 -2 56 2
rect 60 -2 64 2
rect 68 -2 72 2
rect 76 -2 80 2
rect 84 -2 88 2
rect 92 -2 96 2
rect 100 -2 104 2
rect 108 -2 112 2
rect 116 -2 120 2
rect 124 -2 128 2
rect 132 -2 136 2
rect 140 -2 142 2
rect 38 -4 142 -2
<< m2contact >>
rect 64 77 68 81
rect 96 77 100 81
rect 56 70 60 74
rect 72 70 76 74
rect 104 70 108 74
rect 88 63 92 67
rect 80 53 84 57
rect 112 53 116 57
rect 48 43 52 47
rect 72 43 76 47
rect 120 39 124 43
rect 136 42 140 46
rect 56 30 60 34
rect 96 32 100 36
rect 64 24 68 28
rect 104 25 108 29
rect 72 17 76 21
rect 56 10 60 14
rect 64 10 68 14
rect 88 10 92 14
rect 96 10 100 14
rect 120 10 124 14
<< metal2 >>
rect 56 34 60 70
rect 56 14 60 30
rect 64 28 68 77
rect 64 14 68 24
rect 72 47 76 70
rect 72 21 76 43
rect 88 14 92 63
rect 96 36 100 77
rect 96 14 100 32
rect 104 29 108 70
rect 120 14 124 39
rect 56 8 60 10
<< labels >>
rlabel metal1 39 0 39 0 2 Gnd!
rlabel metal1 39 90 39 90 3 Vdd!
rlabel m2contact 138 44 138 44 1 q
rlabel m2contact 50 45 50 45 1 d
rlabel m2contact 74 45 74 45 1 ph2
rlabel m2contact 82 55 82 55 1 ph2b
rlabel m2contact 114 55 114 55 1 ph1b
rlabel m2contact 106 27 106 27 1 ph1
<< end >>
