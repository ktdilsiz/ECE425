magic
tech scmos
timestamp 1484534894
<< metal1 >>
rect -2 856 22 864
rect 8 816 19 820
rect 8 809 12 816
rect -2 766 22 774
rect -2 746 22 754
rect 8 706 19 710
rect 8 699 12 706
rect -2 656 22 664
rect -2 636 22 644
rect 8 596 19 600
rect 8 589 12 596
rect -2 546 22 554
rect -2 526 22 534
rect 8 486 19 490
rect 8 479 12 486
rect -2 436 22 444
rect -2 416 22 424
rect 8 376 19 380
rect 8 369 12 376
rect -2 326 22 334
rect -2 306 22 314
rect 8 266 19 270
rect 8 259 12 266
rect -2 216 22 224
rect -2 196 22 204
rect 8 156 19 160
rect 8 149 12 156
rect -2 106 22 114
rect -2 86 22 94
rect 8 46 19 50
rect 8 39 12 46
rect -2 -4 22 4
<< m2contact >>
rect 0 808 4 812
rect 0 698 4 702
rect 0 588 4 592
rect 0 478 4 482
rect 0 368 4 372
rect 0 258 4 262
rect 0 148 4 152
rect 0 38 4 42
<< metal2 >>
rect -1 842 5 843
rect -1 838 0 842
rect 4 838 5 842
rect -1 837 5 838
rect 47 842 53 843
rect 47 838 48 842
rect 52 838 53 842
rect 47 837 53 838
rect 0 812 4 837
rect 48 815 52 837
rect -1 732 5 733
rect -1 728 0 732
rect 4 728 5 732
rect -1 727 5 728
rect 47 732 53 733
rect 47 728 48 732
rect 52 728 53 732
rect 47 727 53 728
rect 0 702 4 727
rect 48 705 52 727
rect -1 622 5 623
rect -1 618 0 622
rect 4 618 5 622
rect -1 617 5 618
rect 47 622 53 623
rect 47 618 48 622
rect 52 618 53 622
rect 47 617 53 618
rect 0 592 4 617
rect 48 595 52 617
rect -1 512 5 513
rect -1 508 0 512
rect 4 508 5 512
rect -1 507 5 508
rect 47 512 53 513
rect 47 508 48 512
rect 52 508 53 512
rect 47 507 53 508
rect 0 482 4 507
rect 48 485 52 507
rect -1 402 5 403
rect -1 398 0 402
rect 4 398 5 402
rect -1 397 5 398
rect 47 402 53 403
rect 47 398 48 402
rect 52 398 53 402
rect 47 397 53 398
rect 0 372 4 397
rect 48 375 52 397
rect -1 292 5 293
rect -1 288 0 292
rect 4 288 5 292
rect -1 287 5 288
rect 47 292 53 293
rect 47 288 48 292
rect 52 288 53 292
rect 47 287 53 288
rect 0 262 4 287
rect 48 265 52 287
rect -1 182 5 183
rect -1 178 0 182
rect 4 178 5 182
rect -1 177 5 178
rect 47 182 53 183
rect 47 178 48 182
rect 52 178 53 182
rect 47 177 53 178
rect 0 152 4 177
rect 48 155 52 177
rect -1 72 5 73
rect -1 68 0 72
rect 4 68 5 72
rect -1 67 5 68
rect 47 72 53 73
rect 47 68 48 72
rect 52 68 53 72
rect 47 67 53 68
rect 0 42 4 67
rect 48 45 52 67
<< m3contact >>
rect 0 838 4 842
rect 48 838 52 842
rect 0 728 4 732
rect 48 728 52 732
rect 0 618 4 622
rect 48 618 52 622
rect 0 508 4 512
rect 48 508 52 512
rect 0 398 4 402
rect 48 398 52 402
rect 0 288 4 292
rect 48 288 52 292
rect 0 178 4 182
rect 48 178 52 182
rect 0 68 4 72
rect 48 68 52 72
<< metal3 >>
rect -1 842 53 843
rect -1 838 0 842
rect 4 838 48 842
rect 52 838 53 842
rect -1 837 53 838
rect -1 732 53 733
rect -1 728 0 732
rect 4 728 48 732
rect 52 728 53 732
rect -1 727 53 728
rect -1 622 53 623
rect -1 618 0 622
rect 4 618 48 622
rect 52 618 53 622
rect -1 617 53 618
rect -1 512 53 513
rect -1 508 0 512
rect 4 508 48 512
rect 52 508 53 512
rect -1 507 53 508
rect -1 402 53 403
rect -1 398 0 402
rect 4 398 48 402
rect 52 398 53 402
rect -1 397 53 398
rect -1 292 53 293
rect -1 288 0 292
rect 4 288 48 292
rect 52 288 53 292
rect -1 287 53 288
rect -1 182 53 183
rect -1 178 0 182
rect 4 178 48 182
rect 52 178 53 182
rect -1 177 53 178
rect -1 72 53 73
rect -1 68 0 72
rect 4 68 48 72
rect 52 68 53 72
rect -1 67 53 68
use inv_1x_8  inv_1x_8_0
timestamp 1484534894
transform 1 0 0 0 1 0
box -6 -4 18 866
use mux2_1x_8  mux2_1x_8_0
timestamp 1484532969
transform 1 0 16 0 1 0
box -6 -4 50 976
<< end >>
