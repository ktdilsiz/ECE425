magic
tech scmos
timestamp 1487714445
<< nwell >>
rect -6 40 50 96
<< ntransistor >>
rect 5 7 7 19
rect 10 7 12 19
rect 18 7 20 19
rect 37 7 39 34
<< ptransistor >>
rect 5 65 7 83
rect 13 65 15 83
rect 21 65 23 83
rect 37 46 39 83
<< ndiffusion >>
rect 32 32 37 34
rect 0 17 5 19
rect 4 8 5 17
rect 0 7 5 8
rect 7 7 10 19
rect 12 17 18 19
rect 12 8 13 17
rect 17 8 18 17
rect 12 7 18 8
rect 20 17 25 19
rect 20 8 21 17
rect 20 7 25 8
rect 36 8 37 32
rect 32 7 37 8
rect 39 32 44 34
rect 39 8 40 32
rect 39 7 44 8
<< pdiffusion >>
rect 0 81 5 83
rect 4 67 5 81
rect 0 65 5 67
rect 7 81 13 83
rect 7 67 8 81
rect 12 67 13 81
rect 7 65 13 67
rect 15 81 21 83
rect 15 67 16 81
rect 20 67 21 81
rect 15 65 21 67
rect 23 81 28 83
rect 23 67 24 81
rect 23 65 28 67
rect 32 81 37 83
rect 36 47 37 81
rect 32 46 37 47
rect 39 81 44 83
rect 39 48 40 81
rect 39 46 44 48
<< ndcontact >>
rect 0 8 4 17
rect 13 8 17 17
rect 21 8 25 17
rect 32 8 36 32
rect 40 8 44 32
<< pdcontact >>
rect 0 67 4 81
rect 8 67 12 81
rect 16 67 20 81
rect 24 67 28 81
rect 32 47 36 81
rect 40 48 44 81
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
rect 40 -2 44 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
rect 32 88 36 92
rect 40 88 44 92
<< polysilicon >>
rect 5 83 7 85
rect 13 83 15 85
rect 21 83 23 85
rect 37 83 39 85
rect 5 63 7 65
rect 13 63 15 65
rect 21 63 23 65
rect 0 61 7 63
rect 10 61 15 63
rect 18 61 23 63
rect 0 47 2 61
rect 10 47 12 61
rect 18 47 20 61
rect 0 23 2 43
rect 0 21 7 23
rect 5 19 7 21
rect 10 19 12 43
rect 18 19 20 43
rect 37 41 39 46
rect 37 34 39 37
rect 5 5 7 7
rect 10 5 12 7
rect 18 5 20 7
rect 37 5 39 7
<< polycontact >>
rect 0 43 4 47
rect 8 43 12 47
rect 16 43 20 47
rect 35 37 39 41
<< metal1 >>
rect -2 92 46 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 32 92
rect 36 88 40 92
rect 44 88 46 92
rect -2 86 46 88
rect 0 81 4 83
rect 0 62 4 67
rect 8 81 12 86
rect 8 65 12 67
rect 16 81 20 83
rect 16 62 20 67
rect 0 58 20 62
rect 24 81 28 83
rect 24 41 28 67
rect 32 81 36 86
rect 32 46 36 47
rect 40 81 44 83
rect 24 37 35 41
rect 24 26 28 37
rect 13 22 28 26
rect 32 32 36 34
rect 0 17 4 19
rect 0 4 4 8
rect 13 17 17 22
rect 13 7 17 8
rect 21 17 25 19
rect 21 4 25 8
rect 32 4 36 8
rect 40 7 44 8
rect -2 2 46 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 40 2
rect 44 -2 46 2
rect -2 -4 46 -2
<< m2contact >>
rect 0 43 4 47
rect 8 43 12 47
rect 16 43 20 47
rect 40 48 44 50
rect 40 46 44 48
rect 40 32 44 34
rect 40 30 44 32
<< metal2 >>
rect 40 34 44 46
<< labels >>
rlabel m2contact 2 45 2 45 1 a
rlabel m2contact 10 45 10 45 1 b
rlabel m2contact 18 45 18 45 1 c
rlabel m2contact 42 48 42 48 1 y
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel metal1 -1 0 -1 0 3 Gnd!
<< end >>
