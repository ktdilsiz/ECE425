magic
tech scmos
timestamp 1487099595
use mux4_dp_1x  mux4_dp_1x_0
array 0 0 112 0 7 112
timestamp 1484419186
transform 1 0 6 0 1 4
box -6 -4 106 96
<< end >>
