magic
tech scmos
timestamp 1494266977
<< m2contact >>
rect -7 -2 7 2
<< end >>
