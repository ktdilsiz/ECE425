magic
tech scmos
timestamp 1484408212
<< end >>
