magic
tech scmos
timestamp 1494278851
<< metal1 >>
rect 162 348 437 351
rect 30 325 642 340
rect 55 300 617 315
rect 55 287 617 293
rect 459 262 469 265
rect 449 257 454 261
rect 217 251 230 253
rect 346 251 357 254
rect 217 248 237 251
rect 323 244 326 249
rect 546 243 550 252
rect 562 243 566 252
rect 146 228 153 236
rect 223 228 230 236
rect 242 228 249 236
rect 386 232 390 242
rect 410 232 414 242
rect 418 239 429 242
rect 535 228 542 236
rect 298 198 309 201
rect 30 187 642 193
rect 339 178 349 181
rect 130 158 134 168
rect 527 148 541 151
rect 451 142 469 145
rect 527 144 534 148
rect 234 136 245 139
rect 218 128 237 131
rect 322 128 326 137
rect 370 112 374 122
rect 55 87 617 93
rect 55 65 617 80
rect 30 40 642 55
<< metal2 >>
rect 18 377 45 380
rect 18 178 21 377
rect 18 3 21 151
rect 30 40 45 340
rect 55 65 70 315
rect 82 151 85 254
rect 162 247 165 351
rect 170 238 173 254
rect 146 218 149 231
rect 82 148 93 151
rect 90 119 93 148
rect 138 138 141 171
rect 130 128 134 137
rect 154 58 157 201
rect 186 181 189 380
rect 242 278 245 321
rect 258 268 301 271
rect 202 248 206 257
rect 176 178 189 181
rect 194 171 197 211
rect 210 178 213 241
rect 170 168 197 171
rect 162 125 165 151
rect 170 137 173 168
rect 186 118 189 145
rect 202 121 205 151
rect 218 128 221 201
rect 226 128 229 231
rect 234 136 237 251
rect 258 247 261 268
rect 202 118 237 121
rect 242 118 245 231
rect 266 198 269 257
rect 282 178 285 251
rect 290 198 293 254
rect 298 178 301 268
rect 322 246 325 261
rect 322 228 325 241
rect 330 221 333 380
rect 434 278 437 351
rect 482 281 485 380
rect 586 377 629 380
rect 482 278 496 281
rect 338 268 349 271
rect 338 238 341 268
rect 346 251 349 268
rect 330 218 341 221
rect 306 181 309 201
rect 306 178 317 181
rect 306 148 309 171
rect 314 138 317 178
rect 330 148 333 181
rect 18 0 45 3
rect 234 0 237 118
rect 258 108 261 132
rect 266 98 269 124
rect 290 98 293 128
rect 322 98 325 131
rect 338 117 341 218
rect 362 198 365 251
rect 370 228 373 261
rect 378 208 381 243
rect 386 218 389 241
rect 402 201 405 264
rect 450 241 453 261
rect 426 238 453 241
rect 394 198 405 201
rect 394 131 397 198
rect 437 178 440 191
rect 386 128 405 131
rect 338 114 365 117
rect 378 108 381 123
rect 394 98 397 123
rect 426 118 430 126
rect 426 101 429 118
rect 434 108 437 132
rect 450 128 453 238
rect 466 178 469 265
rect 474 218 477 254
rect 482 238 485 251
rect 506 238 509 254
rect 490 208 493 231
rect 514 211 517 254
rect 546 248 549 271
rect 562 248 565 271
rect 586 268 589 377
rect 522 228 525 244
rect 506 208 517 211
rect 474 148 477 201
rect 458 125 461 141
rect 506 121 509 208
rect 538 148 541 231
rect 570 181 573 251
rect 586 188 589 254
rect 570 178 586 181
rect 426 98 437 101
rect 434 0 437 98
rect 570 58 573 112
rect 586 3 589 134
rect 602 65 617 315
rect 627 40 642 340
rect 666 248 669 321
rect 586 0 629 3
<< metal3 >>
rect 0 317 246 322
rect 667 317 672 322
rect 337 267 550 272
rect 561 267 590 272
rect 129 257 326 262
rect 369 257 582 262
rect 201 247 670 252
rect 169 237 214 242
rect 321 237 414 242
rect 481 237 510 242
rect 105 227 526 232
rect 145 217 182 222
rect 337 217 478 222
rect 193 207 382 212
rect 465 207 494 212
rect 217 197 366 202
rect 473 197 529 202
rect 0 187 441 192
rect 585 187 672 192
rect 17 177 254 182
rect 281 177 334 182
rect 345 177 470 182
rect 281 172 286 177
rect 137 167 286 172
rect 305 167 521 172
rect 129 157 542 162
rect 17 147 86 152
rect 121 147 510 152
rect 313 137 462 142
rect 97 127 518 132
rect 185 117 374 122
rect 257 107 590 112
rect 265 97 430 102
rect 0 57 158 62
rect 569 57 672 62
use $$M2_M1  $$M2_M1_0
timestamp 1494266977
transform 1 0 164 0 1 350
box -2 -2 2 2
use $$M2_M1  $$M2_M1_1
timestamp 1494266977
transform 1 0 436 0 1 350
box -2 -2 2 2
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_0
timestamp 1494266977
transform 1 0 37 0 1 332
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_1
timestamp 1494266977
transform 1 0 634 0 1 332
box -7 -7 7 7
use $$M3_M2  $$M3_M2_0
timestamp 1494266977
transform 1 0 244 0 1 320
box -3 -3 3 3
use $$M3_M2  $$M3_M2_1
timestamp 1494266977
transform 1 0 668 0 1 320
box -3 -3 3 3
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_2
timestamp 1494266977
transform 1 0 62 0 1 307
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_3
timestamp 1494266977
transform 1 0 609 0 1 307
box -7 -7 7 7
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_0
timestamp 1494266977
transform 1 0 62 0 1 290
box -7 -2 7 2
use $$M3_M2  $$M3_M2_2
timestamp 1494266977
transform 1 0 132 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_3
timestamp 1494266977
transform 1 0 84 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_2
timestamp 1494266977
transform 1 0 132 0 1 256
box -2 -2 2 2
use $$M2_M1  $$M2_M1_4
timestamp 1494266977
transform 1 0 108 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_3
timestamp 1494266977
transform 1 0 108 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_5
timestamp 1494266977
transform 1 0 172 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_6
timestamp 1494266977
transform 1 0 188 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_7
timestamp 1494266977
transform 1 0 164 0 1 249
box -2 -2 2 2
use $$M2_M1  $$M2_M1_8
timestamp 1494266977
transform 1 0 148 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_5
timestamp 1494266977
transform 1 0 148 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_4
timestamp 1494266977
transform 1 0 172 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_9
timestamp 1494266977
transform 1 0 180 0 1 220
box -2 -2 2 2
use $$M3_M2  $$M3_M2_6
timestamp 1494266977
transform 1 0 180 0 1 220
box -3 -3 3 3
use $$M2_M1  $$M2_M1_10
timestamp 1494266977
transform 1 0 158 0 1 200
box -2 -2 2 2
use $$M2_M1  $$M2_M1_11
timestamp 1494266977
transform 1 0 204 0 1 255
box -2 -2 2 2
use $$M3_M2  $$M3_M2_7
timestamp 1494266977
transform 1 0 204 0 1 250
box -3 -3 3 3
use $$M3_M2  $$M3_M2_10
timestamp 1494266977
transform 1 0 196 0 1 210
box -3 -3 3 3
use $$M2_M1  $$M2_M1_16
timestamp 1494266977
transform 1 0 212 0 1 243
box -2 -2 2 2
use $$M3_M2  $$M3_M2_9
timestamp 1494266977
transform 1 0 212 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_12
timestamp 1494266977
transform 1 0 244 0 1 280
box -2 -2 2 2
use $$M2_M1  $$M2_M1_13
timestamp 1494266977
transform 1 0 236 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_17
timestamp 1494266977
transform 1 0 228 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_11
timestamp 1494266977
transform 1 0 220 0 1 200
box -3 -3 3 3
use $$M2_M1  $$M2_M1_14
timestamp 1494266977
transform 1 0 276 0 1 260
box -2 -2 2 2
use $$M2_M1  $$M2_M1_15
timestamp 1494266977
transform 1 0 268 0 1 256
box -2 -2 2 2
use $$M3_M2  $$M3_M2_8
timestamp 1494266977
transform 1 0 276 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_18
timestamp 1494266977
transform 1 0 260 0 1 249
box -2 -2 2 2
use $$M2_M1  $$M2_M1_19
timestamp 1494266977
transform 1 0 244 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_12
timestamp 1494266977
transform 1 0 268 0 1 200
box -3 -3 3 3
use $$M2_M1  $$M2_M1_20
timestamp 1494266977
transform 1 0 284 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_21
timestamp 1494266977
transform 1 0 292 0 1 253
box -2 -2 2 2
use $$M3_M2  $$M3_M2_13
timestamp 1494266977
transform 1 0 284 0 1 250
box -3 -3 3 3
use $$M3_M2  $$M3_M2_14
timestamp 1494266977
transform 1 0 292 0 1 200
box -3 -3 3 3
use $$M2_M1  $$M2_M1_27
timestamp 1494266977
transform 1 0 308 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_15
timestamp 1494266977
transform 1 0 340 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_16
timestamp 1494266977
transform 1 0 324 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_23
timestamp 1494266977
transform 1 0 324 0 1 248
box -2 -2 2 2
use $$M3_M2  $$M3_M2_17
timestamp 1494266977
transform 1 0 324 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_22
timestamp 1494266977
transform 1 0 348 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_24
timestamp 1494266977
transform 1 0 340 0 1 240
box -2 -2 2 2
use $$M2_M1  $$M2_M1_25
timestamp 1494266977
transform 1 0 324 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_18
timestamp 1494266977
transform 1 0 340 0 1 220
box -3 -3 3 3
use $$M2_M1  $$M2_M1_26
timestamp 1494266977
transform 1 0 332 0 1 210
box -2 -2 2 2
use $$M3_M2  $$M3_M2_19
timestamp 1494266977
transform 1 0 332 0 1 210
box -3 -3 3 3
use $$M3_M2  $$M3_M2_20
timestamp 1494266977
transform 1 0 372 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_28
timestamp 1494266977
transform 1 0 364 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_29
timestamp 1494266977
transform 1 0 380 0 1 241
box -2 -2 2 2
use $$M2_M1  $$M2_M1_30
timestamp 1494266977
transform 1 0 396 0 1 264
box -2 -2 2 2
use $$M3_M2  $$M3_M2_21
timestamp 1494266977
transform 1 0 396 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_31
timestamp 1494266977
transform 1 0 404 0 1 263
box -2 -2 2 2
use $$M2_M1  $$M2_M1_32
timestamp 1494266977
transform 1 0 388 0 1 240
box -2 -2 2 2
use $$M2_M1  $$M2_M1_33
timestamp 1494266977
transform 1 0 372 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_22
timestamp 1494266977
transform 1 0 388 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_23
timestamp 1494266977
transform 1 0 380 0 1 210
box -3 -3 3 3
use $$M3_M2  $$M3_M2_24
timestamp 1494266977
transform 1 0 364 0 1 200
box -3 -3 3 3
use $$M2_M1  $$M2_M1_37
timestamp 1494266977
transform 1 0 412 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_25
timestamp 1494266977
transform 1 0 412 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_34
timestamp 1494266977
transform 1 0 436 0 1 280
box -2 -2 2 2
use $$M2_M1  $$M2_M1_38
timestamp 1494266977
transform 1 0 428 0 1 240
box -2 -2 2 2
use $$M2_M1  $$M2_M1_36
timestamp 1494266977
transform 1 0 452 0 1 260
box -2 -2 2 2
use $$M2_M1  $$M2_M1_35
timestamp 1494266977
transform 1 0 468 0 1 264
box -2 -2 2 2
use $$M2_M1  $$M2_M1_39
timestamp 1494266977
transform 1 0 495 0 1 280
box -2 -2 2 2
use $$M2_M1  $$M2_M1_40
timestamp 1494266977
transform 1 0 476 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_41
timestamp 1494266977
transform 1 0 484 0 1 250
box -2 -2 2 2
use $$M3_M2  $$M3_M2_26
timestamp 1494266977
transform 1 0 484 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_42
timestamp 1494266977
transform 1 0 492 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_27
timestamp 1494266977
transform 1 0 476 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_28
timestamp 1494266977
transform 1 0 468 0 1 210
box -3 -3 3 3
use $$M3_M2  $$M3_M2_29
timestamp 1494266977
transform 1 0 492 0 1 210
box -3 -3 3 3
use $$M3_M2  $$M3_M2_30
timestamp 1494266977
transform 1 0 476 0 1 200
box -3 -3 3 3
use $$M2_M1  $$M2_M1_43
timestamp 1494266977
transform 1 0 508 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_44
timestamp 1494266977
transform 1 0 516 0 1 253
box -2 -2 2 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_1
timestamp 1494266977
transform 1 0 609 0 1 290
box -7 -2 7 2
use $$M3_M2  $$M3_M2_32
timestamp 1494266977
transform 1 0 548 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_33
timestamp 1494266977
transform 1 0 564 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_34
timestamp 1494266977
transform 1 0 588 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_31
timestamp 1494266977
transform 1 0 508 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_45
timestamp 1494266977
transform 1 0 524 0 1 243
box -2 -2 2 2
use $$M3_M2  $$M3_M2_36
timestamp 1494266977
transform 1 0 524 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_46
timestamp 1494266977
transform 1 0 580 0 1 260
box -2 -2 2 2
use $$M3_M2  $$M3_M2_35
timestamp 1494266977
transform 1 0 580 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_48
timestamp 1494266977
transform 1 0 548 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_49
timestamp 1494266977
transform 1 0 564 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_50
timestamp 1494266977
transform 1 0 572 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_47
timestamp 1494266977
transform 1 0 588 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_51
timestamp 1494266977
transform 1 0 540 0 1 230
box -2 -2 2 2
use $$M2_M1  $$M2_M1_52
timestamp 1494266977
transform 1 0 527 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_37
timestamp 1494266977
transform 1 0 527 0 1 200
box -3 -3 3 3
use $$M3_M2  $$M3_M2_38
timestamp 1494266977
transform 1 0 668 0 1 250
box -3 -3 3 3
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_2
timestamp 1494266977
transform 1 0 37 0 1 190
box -7 -2 7 2
use XNOR2X1  XNOR2X1_0
timestamp 1494266853
transform -1 0 136 0 -1 290
box -8 -3 64 105
use FILL  FILL_0
timestamp 1494266977
transform 1 0 136 0 -1 290
box -8 -3 16 105
use OAI21X1  OAI21X1_0
timestamp 1494266977
transform -1 0 176 0 -1 290
box -8 -3 34 105
use INVX2  INVX2_0
timestamp 1494266977
transform -1 0 192 0 -1 290
box -9 -3 26 105
use FILL  FILL_1
timestamp 1494266977
transform 1 0 192 0 -1 290
box -8 -3 16 105
use OAI21X1  OAI21X1_1
timestamp 1494266977
transform 1 0 200 0 -1 290
box -8 -3 34 105
use FILL  FILL_2
timestamp 1494266977
transform 1 0 232 0 -1 290
box -8 -3 16 105
use OAI21X1  OAI21X1_2
timestamp 1494266977
transform -1 0 272 0 -1 290
box -8 -3 34 105
use INVX2  INVX2_1
timestamp 1494266977
transform -1 0 288 0 -1 290
box -9 -3 26 105
use INVX2  INVX2_2
timestamp 1494266977
transform 1 0 288 0 -1 290
box -9 -3 26 105
use FILL  FILL_3
timestamp 1494266977
transform 1 0 304 0 -1 290
box -8 -3 16 105
use NAND3X1  NAND3X1_0
timestamp 1494266977
transform -1 0 344 0 -1 290
box -8 -3 40 105
use FILL  FILL_4
timestamp 1494266977
transform 1 0 344 0 -1 290
box -8 -3 16 105
use NAND2X1  NAND2X1_0
timestamp 1494266977
transform 1 0 352 0 -1 290
box -8 -3 32 105
use NOR2X1  NOR2X1_0
timestamp 1494266977
transform -1 0 400 0 -1 290
box -8 -3 32 105
use NOR2X1  NOR2X1_1
timestamp 1494266977
transform 1 0 400 0 -1 290
box -8 -3 32 105
use $$M3_M2  $$M3_M2_39
timestamp 1494266977
transform 1 0 439 0 1 190
box -3 -3 3 3
use FILL  FILL_5
timestamp 1494266977
transform 1 0 424 0 -1 290
box -8 -3 16 105
use OR2X1  OR2X1_0
timestamp 1494266977
transform -1 0 464 0 -1 290
box -8 -3 40 105
use FILL  FILL_6
timestamp 1494266977
transform 1 0 464 0 -1 290
box -8 -3 16 105
use INVX2  INVX2_3
timestamp 1494266977
transform 1 0 472 0 -1 290
box -9 -3 26 105
use NAND2X1  NAND2X1_1
timestamp 1494266977
transform -1 0 512 0 -1 290
box -8 -3 32 105
use OAI21X1  OAI21X1_3
timestamp 1494266977
transform 1 0 512 0 -1 290
box -8 -3 34 105
use AND2X2  AND2X2_0
timestamp 1494266977
transform -1 0 576 0 -1 290
box -8 -3 40 105
use $$M3_M2  $$M3_M2_40
timestamp 1494266977
transform 1 0 588 0 1 190
box -3 -3 3 3
use INVX2  INVX2_4
timestamp 1494266977
transform -1 0 592 0 -1 290
box -9 -3 26 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_3
timestamp 1494266977
transform 1 0 634 0 1 190
box -7 -2 7 2
use $$M3_M2  $$M3_M2_41
timestamp 1494266977
transform 1 0 20 0 1 180
box -3 -3 3 3
use $$M3_M2  $$M3_M2_42
timestamp 1494266977
transform 1 0 20 0 1 150
box -3 -3 3 3
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_4
timestamp 1494266977
transform 1 0 62 0 1 90
box -7 -2 7 2
use $$M3_M2  $$M3_M2_43
timestamp 1494266977
transform 1 0 84 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_53
timestamp 1494266977
transform 1 0 100 0 1 130
box -2 -2 2 2
use $$M3_M2  $$M3_M2_44
timestamp 1494266977
transform 1 0 100 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_54
timestamp 1494266977
transform 1 0 92 0 1 121
box -2 -2 2 2
use FILL  FILL_7
timestamp 1494266977
transform -1 0 88 0 1 90
box -8 -3 16 105
use INVX2  INVX2_5
timestamp 1494266977
transform 1 0 88 0 1 90
box -9 -3 26 105
use FILL  FILL_8
timestamp 1494266977
transform -1 0 112 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_45
timestamp 1494266977
transform 1 0 140 0 1 170
box -3 -3 3 3
use $$M2_M1  $$M2_M1_56
timestamp 1494266977
transform 1 0 132 0 1 160
box -2 -2 2 2
use $$M3_M2  $$M3_M2_46
timestamp 1494266977
transform 1 0 132 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_57
timestamp 1494266977
transform 1 0 124 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_47
timestamp 1494266977
transform 1 0 124 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_59
timestamp 1494266977
transform 1 0 140 0 1 140
box -2 -2 2 2
use $$M2_M1  $$M2_M1_61
timestamp 1494266977
transform 1 0 132 0 1 135
box -2 -2 2 2
use $$M3_M2  $$M3_M2_49
timestamp 1494266977
transform 1 0 132 0 1 130
box -3 -3 3 3
use NAND3X1  NAND3X1_1
timestamp 1494266977
transform -1 0 144 0 1 90
box -8 -3 40 105
use FILL  FILL_9
timestamp 1494266977
transform -1 0 152 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_55
timestamp 1494266977
transform 1 0 177 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_48
timestamp 1494266977
transform 1 0 164 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_58
timestamp 1494266977
transform 1 0 188 0 1 144
box -2 -2 2 2
use $$M2_M1  $$M2_M1_60
timestamp 1494266977
transform 1 0 172 0 1 139
box -2 -2 2 2
use $$M2_M1  $$M2_M1_62
timestamp 1494266977
transform 1 0 164 0 1 127
box -2 -2 2 2
use FILL  FILL_10
timestamp 1494266977
transform -1 0 160 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_50
timestamp 1494266977
transform 1 0 188 0 1 120
box -3 -3 3 3
use OAI21X1  OAI21X1_4
timestamp 1494266977
transform 1 0 160 0 1 90
box -8 -3 34 105
use $$M2_M1  $$M2_M1_63
timestamp 1494266977
transform 1 0 212 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_53
timestamp 1494266977
transform 1 0 204 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_75
timestamp 1494266977
transform 1 0 204 0 1 121
box -2 -2 2 2
use FILL  FILL_11
timestamp 1494266977
transform -1 0 200 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_64
timestamp 1494266977
transform 1 0 252 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_51
timestamp 1494266977
transform 1 0 252 0 1 180
box -3 -3 3 3
use $$M2_M1  $$M2_M1_66
timestamp 1494266977
transform 1 0 236 0 1 137
box -2 -2 2 2
use $$M2_M1  $$M2_M1_68
timestamp 1494266977
transform 1 0 220 0 1 130
box -2 -2 2 2
use $$M3_M2  $$M3_M2_54
timestamp 1494266977
transform 1 0 228 0 1 130
box -3 -3 3 3
use INVX2  INVX2_6
timestamp 1494266977
transform 1 0 200 0 1 90
box -9 -3 26 105
use FILL  FILL_12
timestamp 1494266977
transform -1 0 224 0 1 90
box -8 -3 16 105
use FILL  FILL_13
timestamp 1494266977
transform -1 0 232 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_67
timestamp 1494266977
transform 1 0 260 0 1 131
box -2 -2 2 2
use $$M3_M2  $$M3_M2_59
timestamp 1494266977
transform 1 0 244 0 1 120
box -3 -3 3 3
use $$M2_M1  $$M2_M1_74
timestamp 1494266977
transform 1 0 268 0 1 123
box -2 -2 2 2
use $$M3_M2  $$M3_M2_60
timestamp 1494266977
transform 1 0 260 0 1 110
box -3 -3 3 3
use $$M3_M2  $$M3_M2_61
timestamp 1494266977
transform 1 0 268 0 1 100
box -3 -3 3 3
use OAI22X1  OAI22X1_0
timestamp 1494266853
transform -1 0 272 0 1 90
box -8 -3 46 105
use $$M3_M2  $$M3_M2_52
timestamp 1494266977
transform 1 0 284 0 1 180
box -3 -3 3 3
use FILL  FILL_14
timestamp 1494266977
transform -1 0 280 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_65
timestamp 1494266977
transform 1 0 300 0 1 180
box -2 -2 2 2
use $$M2_M1  $$M2_M1_73
timestamp 1494266977
transform 1 0 292 0 1 127
box -2 -2 2 2
use $$M3_M2  $$M3_M2_62
timestamp 1494266977
transform 1 0 292 0 1 100
box -3 -3 3 3
use FILL  FILL_15
timestamp 1494266977
transform -1 0 288 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_55
timestamp 1494266977
transform 1 0 332 0 1 180
box -3 -3 3 3
use $$M3_M2  $$M3_M2_57
timestamp 1494266977
transform 1 0 308 0 1 170
box -3 -3 3 3
use $$M2_M1  $$M2_M1_70
timestamp 1494266977
transform 1 0 308 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_71
timestamp 1494266977
transform 1 0 332 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_72
timestamp 1494266977
transform 1 0 316 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_58
timestamp 1494266977
transform 1 0 316 0 1 140
box -3 -3 3 3
use NAND2X1  NAND2X1_2
timestamp 1494266977
transform 1 0 288 0 1 90
box -8 -3 32 105
use $$M2_M1  $$M2_M1_76
timestamp 1494266977
transform 1 0 324 0 1 130
box -2 -2 2 2
use $$M3_M2  $$M3_M2_63
timestamp 1494266977
transform 1 0 324 0 1 100
box -3 -3 3 3
use $$M2_M1  $$M2_M1_69
timestamp 1494266977
transform 1 0 348 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_56
timestamp 1494266977
transform 1 0 348 0 1 180
box -3 -3 3 3
use NAND3X1  NAND3X1_2
timestamp 1494266977
transform 1 0 312 0 1 90
box -8 -3 40 105
use FILL  FILL_16
timestamp 1494266977
transform -1 0 352 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_77
timestamp 1494266977
transform 1 0 388 0 1 133
box -2 -2 2 2
use $$M2_M1  $$M2_M1_81
timestamp 1494266977
transform 1 0 372 0 1 120
box -2 -2 2 2
use $$M2_M1  $$M2_M1_78
timestamp 1494266977
transform 1 0 380 0 1 122
box -2 -2 2 2
use $$M3_M2  $$M3_M2_64
timestamp 1494266977
transform 1 0 372 0 1 120
box -3 -3 3 3
use $$M2_M1  $$M2_M1_80
timestamp 1494266977
transform 1 0 396 0 1 121
box -2 -2 2 2
use $$M2_M1  $$M2_M1_82
timestamp 1494266977
transform 1 0 364 0 1 115
box -2 -2 2 2
use FILL  FILL_17
timestamp 1494266977
transform -1 0 360 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_65
timestamp 1494266977
transform 1 0 380 0 1 110
box -3 -3 3 3
use $$M3_M2  $$M3_M2_66
timestamp 1494266977
transform 1 0 396 0 1 100
box -3 -3 3 3
use AOI21X1  AOI21X1_0
timestamp 1494266977
transform -1 0 392 0 1 90
box -7 -3 39 105
use $$M2_M1  $$M2_M1_79
timestamp 1494266977
transform 1 0 404 0 1 130
box -2 -2 2 2
use INVX2  INVX2_7
timestamp 1494266977
transform 1 0 392 0 1 90
box -9 -3 26 105
use FILL  FILL_18
timestamp 1494266977
transform -1 0 416 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_83
timestamp 1494266977
transform 1 0 439 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_67
timestamp 1494266977
transform 1 0 468 0 1 180
box -3 -3 3 3
use $$M2_M1  $$M2_M1_85
timestamp 1494266977
transform 1 0 476 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_68
timestamp 1494266977
transform 1 0 460 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_84
timestamp 1494266977
transform 1 0 436 0 1 131
box -2 -2 2 2
use $$M2_M1  $$M2_M1_86
timestamp 1494266977
transform 1 0 428 0 1 124
box -2 -2 2 2
use $$M3_M2  $$M3_M2_69
timestamp 1494266977
transform 1 0 452 0 1 130
box -3 -3 3 3
use $$M3_M2  $$M3_M2_70
timestamp 1494266977
transform 1 0 436 0 1 110
box -3 -3 3 3
use $$M3_M2  $$M3_M2_71
timestamp 1494266977
transform 1 0 428 0 1 100
box -3 -3 3 3
use FILL  FILL_19
timestamp 1494266977
transform -1 0 424 0 1 90
box -8 -3 16 105
use OAI21X1  OAI21X1_5
timestamp 1494266977
transform 1 0 424 0 1 90
box -8 -3 34 105
use $$M2_M1  $$M2_M1_87
timestamp 1494266977
transform 1 0 460 0 1 127
box -2 -2 2 2
use NAND2X1  NAND2X1_3
timestamp 1494266977
transform 1 0 456 0 1 90
box -8 -3 32 105
use FILL  FILL_20
timestamp 1494266977
transform -1 0 488 0 1 90
box -8 -3 16 105
use FILL  FILL_21
timestamp 1494266977
transform -1 0 496 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_88
timestamp 1494266977
transform 1 0 519 0 1 170
box -2 -2 2 2
use $$M3_M2  $$M3_M2_72
timestamp 1494266977
transform 1 0 519 0 1 170
box -3 -3 3 3
use $$M3_M2  $$M3_M2_74
timestamp 1494266977
transform 1 0 508 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_91
timestamp 1494266977
transform 1 0 516 0 1 131
box -2 -2 2 2
use $$M3_M2  $$M3_M2_75
timestamp 1494266977
transform 1 0 516 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_92
timestamp 1494266977
transform 1 0 508 0 1 123
box -2 -2 2 2
use FILL  FILL_22
timestamp 1494266977
transform -1 0 504 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_73
timestamp 1494266977
transform 1 0 540 0 1 160
box -3 -3 3 3
use OAI21X1  OAI21X1_6
timestamp 1494266977
transform 1 0 504 0 1 90
box -8 -3 34 105
use $$M2_M1  $$M2_M1_90
timestamp 1494266977
transform 1 0 540 0 1 150
box -2 -2 2 2
use FILL  FILL_23
timestamp 1494266977
transform -1 0 544 0 1 90
box -8 -3 16 105
use FILL  FILL_24
timestamp 1494266977
transform -1 0 552 0 1 90
box -8 -3 16 105
use FILL  FILL_25
timestamp 1494266977
transform -1 0 560 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_89
timestamp 1494266977
transform 1 0 585 0 1 180
box -2 -2 2 2
use $$M2_M1  $$M2_M1_93
timestamp 1494266977
transform 1 0 588 0 1 133
box -2 -2 2 2
use $$M2_M1  $$M2_M1_94
timestamp 1494266977
transform 1 0 572 0 1 111
box -2 -2 2 2
use FILL  FILL_26
timestamp 1494266977
transform -1 0 568 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_76
timestamp 1494266977
transform 1 0 588 0 1 110
box -3 -3 3 3
use NOR2X1  NOR2X1_2
timestamp 1494266977
transform 1 0 568 0 1 90
box -8 -3 32 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_5
timestamp 1494266977
transform 1 0 609 0 1 90
box -7 -2 7 2
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_4
timestamp 1494266977
transform 1 0 62 0 1 72
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_5
timestamp 1494266977
transform 1 0 609 0 1 72
box -7 -7 7 7
use $$M3_M2  $$M3_M2_77
timestamp 1494266977
transform 1 0 156 0 1 60
box -3 -3 3 3
use $$M3_M2  $$M3_M2_78
timestamp 1494266977
transform 1 0 572 0 1 60
box -3 -3 3 3
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_6
timestamp 1494266977
transform 1 0 37 0 1 47
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_7
timestamp 1494266977
transform 1 0 634 0 1 47
box -7 -7 7 7
<< labels >>
flabel metal3 2 320 2 320 4 FreeSans 26 0 0 0 alucontrol[4]
flabel metal3 2 190 2 190 4 FreeSans 26 0 0 0 alucontrol[5]
flabel metal3 2 60 2 60 4 FreeSans 26 0 0 0 alucontrol[6]
flabel metal2 332 378 332 378 4 FreeSans 26 0 0 0 alucontrol[1]
flabel metal2 188 378 188 378 4 FreeSans 26 0 0 0 alucontrol[2]
flabel metal2 484 378 484 378 4 FreeSans 26 0 0 0 alucontrol[0]
flabel metal2 44 378 44 378 4 FreeSans 26 0 0 0 alucontrol[3]
flabel metal2 628 378 628 378 4 FreeSans 26 0 0 0 funct[5]
flabel metal3 669 320 669 320 4 FreeSans 26 0 0 0 funct[2]
flabel metal3 669 60 669 60 4 FreeSans 26 0 0 0 funct[4]
flabel metal3 669 190 669 190 4 FreeSans 26 0 0 0 funct[3]
flabel metal2 628 1 628 1 4 FreeSans 26 0 0 0 aluop[0]
flabel metal2 44 1 44 1 4 FreeSans 26 0 0 0 funct[1]
flabel metal2 236 1 236 1 4 FreeSans 26 0 0 0 funct[0]
flabel metal2 436 1 436 1 4 FreeSans 26 0 0 0 aluop[1]
rlabel metal1 263 332 263 332 1 Vdd!
rlabel metal1 266 307 266 307 1 Gnd!
<< end >>
