magic
tech scmos
timestamp 1490727624
<< metal1 >>
rect 30 525 1042 540
rect 55 500 1017 515
rect 55 487 1017 493
rect 106 458 110 467
rect 282 453 286 462
rect 626 453 630 462
rect 790 454 798 462
rect 482 448 493 451
rect 498 443 502 452
rect 514 443 518 452
rect 642 444 677 447
rect 690 443 694 452
rect 699 448 709 451
rect 898 448 903 457
rect 143 428 150 436
rect 410 434 414 442
rect 906 440 933 443
rect 890 428 897 436
rect 210 398 221 401
rect 30 387 1042 393
rect 274 378 283 382
rect 362 378 381 381
rect 890 378 933 381
rect 114 348 125 351
rect 202 348 213 351
rect 210 345 213 348
rect 283 331 293 334
rect 394 328 398 337
rect 442 333 446 342
rect 546 333 581 336
rect 594 328 598 337
rect 730 333 734 342
rect 138 321 149 324
rect 187 321 195 327
rect 178 318 195 321
rect 426 319 431 323
rect 530 318 534 327
rect 634 323 638 332
rect 946 328 950 337
rect 650 321 665 324
rect 682 321 686 327
rect 690 323 709 326
rect 690 321 693 323
rect 682 318 693 321
rect 745 319 750 323
rect 682 312 686 318
rect 458 308 469 311
rect 55 287 1017 293
rect 754 278 789 281
rect 931 278 949 281
rect 194 268 198 278
rect 282 255 293 258
rect 410 254 418 262
rect 970 258 974 267
rect 115 251 142 254
rect 530 251 534 254
rect 530 248 566 251
rect 746 248 750 257
rect 826 251 829 256
rect 810 248 829 251
rect 841 251 854 253
rect 841 248 861 251
rect 866 248 879 253
rect 891 251 901 254
rect 234 241 245 244
rect 554 243 566 248
rect 659 244 677 247
rect 220 228 225 236
rect 322 232 326 242
rect 666 238 669 241
rect 674 238 677 244
rect 707 238 725 241
rect 490 228 494 237
rect 666 231 670 234
rect 682 231 686 237
rect 514 228 525 231
rect 666 228 686 231
rect 722 231 725 238
rect 722 228 733 231
rect 866 228 873 236
rect 927 228 934 236
rect 30 187 1042 193
rect 237 178 246 182
rect 114 138 118 148
rect 331 142 341 145
rect 348 144 353 152
rect 242 118 246 127
rect 321 123 326 132
rect 338 131 341 142
rect 578 138 582 147
rect 762 144 769 152
rect 610 138 621 141
rect 866 138 870 147
rect 338 128 359 131
rect 346 126 359 128
rect 553 128 573 131
rect 650 128 661 131
rect 553 126 566 128
rect 747 125 757 128
rect 730 121 741 124
rect 394 102 398 112
rect 403 109 413 112
rect 690 102 694 112
rect 410 98 421 101
rect 55 87 1017 93
rect 55 65 1017 80
rect 30 40 1042 55
<< metal2 >>
rect 18 577 45 580
rect 18 478 21 577
rect 2 58 5 161
rect 18 3 21 201
rect 30 40 45 540
rect 55 65 70 515
rect 146 478 149 521
rect 186 478 189 580
rect 90 378 93 401
rect 82 318 93 321
rect 90 257 93 318
rect 106 278 109 461
rect 114 328 117 351
rect 106 198 109 211
rect 114 138 117 161
rect 122 131 125 454
rect 130 378 133 441
rect 178 388 181 454
rect 162 331 165 340
rect 154 328 165 331
rect 146 228 149 324
rect 154 242 157 328
rect 194 311 197 351
rect 202 348 205 361
rect 202 333 206 342
rect 210 328 213 401
rect 194 308 205 311
rect 162 218 165 241
rect 170 208 173 291
rect 202 248 205 308
rect 218 278 221 391
rect 274 378 277 451
rect 282 438 285 461
rect 322 448 325 580
rect 298 378 301 447
rect 330 381 333 521
rect 466 468 469 580
rect 538 457 541 471
rect 602 458 605 580
rect 746 577 749 580
rect 882 577 885 580
rect 986 577 1029 580
rect 320 378 333 381
rect 226 325 229 361
rect 330 342 334 352
rect 242 325 245 341
rect 242 254 245 271
rect 18 0 45 3
rect 186 0 189 211
rect 202 168 205 241
rect 234 131 237 251
rect 242 178 245 244
rect 250 231 253 301
rect 266 261 269 281
rect 266 258 285 261
rect 250 228 261 231
rect 250 114 253 228
rect 266 198 269 258
rect 266 125 269 171
rect 282 148 285 171
rect 218 98 221 111
rect 290 108 293 334
rect 306 325 309 341
rect 378 338 381 401
rect 314 308 317 332
rect 346 319 349 331
rect 298 278 301 301
rect 354 298 357 311
rect 314 218 317 242
rect 354 228 357 264
rect 370 228 373 311
rect 402 278 405 331
rect 418 311 421 321
rect 426 318 429 341
rect 442 338 445 351
rect 418 308 429 311
rect 458 308 461 321
rect 386 228 389 260
rect 410 248 413 261
rect 306 121 309 141
rect 314 135 317 191
rect 346 168 349 201
rect 378 191 381 201
rect 378 188 389 191
rect 322 128 325 161
rect 386 137 389 188
rect 410 158 413 241
rect 322 0 325 121
rect 362 101 365 132
rect 418 128 421 144
rect 426 138 429 308
rect 482 278 485 451
rect 498 418 501 451
rect 666 441 669 451
rect 522 438 533 441
rect 658 438 669 441
rect 522 418 525 438
rect 530 318 533 431
rect 498 248 502 257
rect 490 228 517 231
rect 370 108 373 126
rect 362 98 413 101
rect 442 98 445 124
rect 466 121 469 141
rect 546 135 549 361
rect 562 318 565 341
rect 594 328 597 411
rect 602 328 605 371
rect 554 168 557 264
rect 570 249 573 271
rect 570 241 581 244
rect 562 145 565 181
rect 570 128 573 241
rect 610 228 613 341
rect 642 331 645 401
rect 642 318 653 321
rect 474 98 477 121
rect 466 0 469 91
rect 498 88 501 122
rect 522 98 525 122
rect 538 98 541 124
rect 578 98 581 141
rect 586 108 589 151
rect 594 118 597 221
rect 626 218 629 242
rect 642 178 645 318
rect 650 228 653 271
rect 658 198 661 438
rect 690 408 693 451
rect 746 448 750 457
rect 794 448 797 461
rect 714 378 717 411
rect 738 408 741 441
rect 898 438 901 451
rect 762 368 765 401
rect 890 378 893 431
rect 666 329 669 341
rect 679 328 682 345
rect 746 261 749 321
rect 754 315 757 331
rect 786 328 789 341
rect 794 281 797 351
rect 810 328 813 341
rect 786 278 797 281
rect 818 278 821 361
rect 826 298 829 351
rect 858 318 861 334
rect 794 271 797 278
rect 794 268 837 271
rect 738 258 749 261
rect 738 251 741 258
rect 802 251 806 256
rect 674 178 677 241
rect 602 0 605 141
rect 626 132 630 142
rect 634 118 637 151
rect 698 148 701 244
rect 706 141 709 251
rect 746 231 749 251
rect 738 228 749 231
rect 802 248 813 251
rect 802 221 805 248
rect 834 247 837 268
rect 746 218 805 221
rect 746 151 749 218
rect 850 208 853 234
rect 858 231 861 251
rect 866 238 869 251
rect 874 248 877 351
rect 914 278 917 454
rect 986 451 989 577
rect 938 448 989 451
rect 922 271 925 401
rect 938 368 941 448
rect 954 311 957 331
rect 946 308 957 311
rect 946 278 949 308
rect 922 268 933 271
rect 882 247 885 261
rect 858 228 869 231
rect 794 198 845 201
rect 714 148 749 151
rect 650 128 653 141
rect 698 138 709 141
rect 698 131 701 138
rect 666 88 669 128
rect 746 0 749 148
rect 754 98 757 128
rect 762 108 765 151
rect 778 128 781 138
rect 786 121 789 151
rect 802 138 805 191
rect 818 148 821 181
rect 810 108 813 136
rect 842 128 845 198
rect 850 108 853 161
rect 858 128 861 151
rect 890 138 893 151
rect 882 0 885 121
rect 898 88 901 254
rect 906 231 909 257
rect 906 228 917 231
rect 930 228 933 268
rect 970 258 973 281
rect 914 178 917 228
rect 957 198 973 201
rect 906 138 909 151
rect 914 135 917 161
rect 922 128 925 151
rect 962 118 965 134
rect 946 88 949 118
rect 970 58 973 198
rect 986 3 989 121
rect 1002 65 1017 515
rect 1027 40 1042 540
rect 986 0 1029 3
<< metal3 >>
rect 0 517 150 522
rect 329 517 1072 522
rect 17 477 102 482
rect 169 477 190 482
rect 465 467 542 472
rect 601 457 630 462
rect 601 452 606 457
rect 105 447 134 452
rect 193 447 326 452
rect 456 447 518 452
rect 537 447 606 452
rect 665 447 798 452
rect 537 443 542 447
rect 529 442 542 443
rect 89 437 134 442
rect 281 437 542 442
rect 793 437 902 442
rect 145 427 190 432
rect 529 427 534 437
rect 497 417 678 422
rect 673 412 678 417
rect 593 407 694 412
rect 713 407 742 412
rect 0 397 94 402
rect 561 397 646 402
rect 921 397 1072 402
rect 177 387 222 392
rect 297 377 366 382
rect 601 367 766 372
rect 860 367 942 372
rect 158 357 230 362
rect 545 357 822 362
rect 97 347 878 352
rect 201 337 566 342
rect 609 337 646 342
rect 665 337 734 342
rect 113 327 350 332
rect 393 327 598 332
rect 633 327 683 332
rect 753 327 814 332
rect 833 327 950 332
rect 89 317 182 322
rect 417 317 462 322
rect 561 317 630 322
rect 777 317 862 322
rect 777 312 782 317
rect 233 307 318 312
rect 353 307 782 312
rect 297 297 830 302
rect 0 287 1072 292
rect 105 277 270 282
rect 401 277 446 282
rect 457 277 486 282
rect 817 277 974 282
rect 193 267 926 272
rect 185 257 270 262
rect 329 257 382 262
rect 881 257 974 262
rect 201 247 278 252
rect 409 247 662 252
rect 705 247 742 252
rect 873 247 958 252
rect 153 237 206 242
rect 321 237 558 242
rect 865 237 918 242
rect 145 227 614 232
rect 689 227 742 232
rect 737 222 742 227
rect 161 217 246 222
rect 289 217 318 222
rect 593 217 742 222
rect 105 207 190 212
rect 622 207 806 212
rect 849 207 902 212
rect 17 197 86 202
rect 313 187 382 192
rect 801 187 806 207
rect 521 177 550 182
rect 561 177 776 182
rect 817 177 963 182
rect 521 172 526 177
rect 0 167 6 172
rect 201 167 270 172
rect 281 167 526 172
rect 553 167 1072 172
rect 1 162 6 167
rect 1 157 118 162
rect 321 157 414 162
rect 505 157 918 162
rect 249 147 352 152
rect 481 147 910 152
rect 233 137 614 142
rect 625 137 654 142
rect 705 137 870 142
rect 121 127 422 132
rect 433 127 726 132
rect 777 127 846 132
rect 857 127 982 132
rect 209 117 246 122
rect 321 117 598 122
rect 633 117 886 122
rect 961 117 990 122
rect 105 107 294 112
rect 369 107 398 112
rect 409 107 518 112
rect 585 107 694 112
rect 737 107 766 112
rect 809 107 854 112
rect 441 97 478 102
rect 521 97 582 102
rect 753 97 822 102
rect 465 87 502 92
rect 601 87 950 92
rect 0 57 5 62
rect 969 57 1072 62
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_0
timestamp 1490727624
transform 1 0 37 0 1 532
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_1
timestamp 1490727624
transform 1 0 1034 0 1 532
box -7 -7 7 7
use $$M3_M2  $$M3_M2_0
timestamp 1490727624
transform 1 0 148 0 1 520
box -3 -3 3 3
use $$M3_M2  $$M3_M2_1
timestamp 1490727624
transform 1 0 332 0 1 520
box -3 -3 3 3
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_2
timestamp 1490727624
transform 1 0 62 0 1 507
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_3
timestamp 1490727624
transform 1 0 1009 0 1 507
box -7 -7 7 7
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_0
timestamp 1490727624
transform 1 0 62 0 1 490
box -7 -2 7 2
use $$M3_M2  $$M3_M2_2
timestamp 1490727624
transform 1 0 20 0 1 480
box -3 -3 3 3
use $$M2_M1  $$M2_M1_0
timestamp 1490727624
transform 1 0 100 0 1 480
box -2 -2 2 2
use $$M3_M2  $$M3_M2_3
timestamp 1490727624
transform 1 0 100 0 1 480
box -3 -3 3 3
use $$M2_M1  $$M2_M1_2
timestamp 1490727624
transform 1 0 92 0 1 441
box -2 -2 2 2
use $$M3_M2  $$M3_M2_5
timestamp 1490727624
transform 1 0 92 0 1 440
box -3 -3 3 3
use $$M3_M2  $$M3_M2_6
timestamp 1490727624
transform 1 0 92 0 1 400
box -3 -3 3 3
use $$M2_M1  $$M2_M1_1
timestamp 1490727624
transform 1 0 108 0 1 460
box -2 -2 2 2
use $$M3_M2  $$M3_M2_4
timestamp 1490727624
transform 1 0 108 0 1 450
box -3 -3 3 3
use $$M2_M1  $$M2_M1_4
timestamp 1490727624
transform 1 0 124 0 1 453
box -2 -2 2 2
use $$M2_M1  $$M2_M1_3
timestamp 1490727624
transform 1 0 148 0 1 480
box -2 -2 2 2
use $$M2_M1  $$M2_M1_5
timestamp 1490727624
transform 1 0 132 0 1 449
box -2 -2 2 2
use $$M3_M2  $$M3_M2_7
timestamp 1490727624
transform 1 0 132 0 1 450
box -3 -3 3 3
use $$M3_M2  $$M3_M2_8
timestamp 1490727624
transform 1 0 132 0 1 440
box -3 -3 3 3
use $$M2_M1  $$M2_M1_6
timestamp 1490727624
transform 1 0 148 0 1 430
box -2 -2 2 2
use $$M3_M2  $$M3_M2_9
timestamp 1490727624
transform 1 0 148 0 1 430
box -3 -3 3 3
use $$M2_M1  $$M2_M1_7
timestamp 1490727624
transform 1 0 172 0 1 480
box -2 -2 2 2
use $$M3_M2  $$M3_M2_10
timestamp 1490727624
transform 1 0 172 0 1 480
box -3 -3 3 3
use $$M3_M2  $$M3_M2_11
timestamp 1490727624
transform 1 0 188 0 1 480
box -3 -3 3 3
use $$M2_M1  $$M2_M1_8
timestamp 1490727624
transform 1 0 180 0 1 453
box -2 -2 2 2
use $$M2_M1  $$M2_M1_10
timestamp 1490727624
transform 1 0 188 0 1 430
box -2 -2 2 2
use $$M3_M2  $$M3_M2_13
timestamp 1490727624
transform 1 0 188 0 1 430
box -3 -3 3 3
use $$M2_M1  $$M2_M1_9
timestamp 1490727624
transform 1 0 196 0 1 453
box -2 -2 2 2
use $$M3_M2  $$M3_M2_12
timestamp 1490727624
transform 1 0 196 0 1 450
box -3 -3 3 3
use $$M2_M1  $$M2_M1_16
timestamp 1490727624
transform 1 0 212 0 1 400
box -2 -2 2 2
use $$M2_M1  $$M2_M1_11
timestamp 1490727624
transform 1 0 284 0 1 460
box -2 -2 2 2
use $$M3_M2  $$M3_M2_15
timestamp 1490727624
transform 1 0 276 0 1 450
box -3 -3 3 3
use $$M2_M1  $$M2_M1_15
timestamp 1490727624
transform 1 0 300 0 1 446
box -2 -2 2 2
use $$M3_M2  $$M3_M2_19
timestamp 1490727624
transform 1 0 284 0 1 440
box -3 -3 3 3
use $$M3_M2  $$M3_M2_16
timestamp 1490727624
transform 1 0 324 0 1 450
box -3 -3 3 3
use $$M3_M2  $$M3_M2_14
timestamp 1490727624
transform 1 0 468 0 1 470
box -3 -3 3 3
use $$M3_M2  $$M3_M2_17
timestamp 1490727624
transform 1 0 459 0 1 450
box -3 -3 3 3
use $$M2_M1  $$M2_M1_17
timestamp 1490727624
transform 1 0 459 0 1 447
box -2 -2 2 2
use $$M2_M1  $$M2_M1_18
timestamp 1490727624
transform 1 0 412 0 1 440
box -2 -2 2 2
use $$M3_M2  $$M3_M2_20
timestamp 1490727624
transform 1 0 412 0 1 440
box -3 -3 3 3
use $$M2_M1  $$M2_M1_21
timestamp 1490727624
transform 1 0 380 0 1 400
box -2 -2 2 2
use $$M2_M1  $$M2_M1_12
timestamp 1490727624
transform 1 0 484 0 1 450
box -2 -2 2 2
use $$M2_M1  $$M2_M1_13
timestamp 1490727624
transform 1 0 500 0 1 450
box -2 -2 2 2
use $$M2_M1  $$M2_M1_14
timestamp 1490727624
transform 1 0 516 0 1 450
box -2 -2 2 2
use $$M3_M2  $$M3_M2_18
timestamp 1490727624
transform 1 0 516 0 1 450
box -3 -3 3 3
use $$M3_M2  $$M3_M2_23
timestamp 1490727624
transform 1 0 500 0 1 420
box -3 -3 3 3
use $$M3_M2  $$M3_M2_21
timestamp 1490727624
transform 1 0 540 0 1 470
box -3 -3 3 3
use $$M2_M1  $$M2_M1_19
timestamp 1490727624
transform 1 0 540 0 1 459
box -2 -2 2 2
use $$M2_M1  $$M2_M1_20
timestamp 1490727624
transform 1 0 532 0 1 440
box -2 -2 2 2
use $$M3_M2  $$M3_M2_22
timestamp 1490727624
transform 1 0 532 0 1 430
box -3 -3 3 3
use $$M3_M2  $$M3_M2_24
timestamp 1490727624
transform 1 0 524 0 1 420
box -3 -3 3 3
use $$M3_M2  $$M3_M2_25
timestamp 1490727624
transform 1 0 604 0 1 460
box -3 -3 3 3
use $$M2_M1  $$M2_M1_22
timestamp 1490727624
transform 1 0 628 0 1 460
box -2 -2 2 2
use $$M3_M2  $$M3_M2_26
timestamp 1490727624
transform 1 0 628 0 1 460
box -3 -3 3 3
use $$M3_M2  $$M3_M2_28
timestamp 1490727624
transform 1 0 596 0 1 410
box -3 -3 3 3
use $$M2_M1  $$M2_M1_24
timestamp 1490727624
transform 1 0 564 0 1 400
box -2 -2 2 2
use $$M3_M2  $$M3_M2_30
timestamp 1490727624
transform 1 0 564 0 1 400
box -3 -3 3 3
use $$M3_M2  $$M3_M2_31
timestamp 1490727624
transform 1 0 644 0 1 400
box -3 -3 3 3
use $$M3_M2  $$M3_M2_27
timestamp 1490727624
transform 1 0 668 0 1 450
box -3 -3 3 3
use $$M2_M1  $$M2_M1_23
timestamp 1490727624
transform 1 0 692 0 1 450
box -2 -2 2 2
use $$M3_M2  $$M3_M2_29
timestamp 1490727624
transform 1 0 692 0 1 410
box -3 -3 3 3
use $$M2_M1  $$M2_M1_25
timestamp 1490727624
transform 1 0 748 0 1 455
box -2 -2 2 2
use $$M3_M2  $$M3_M2_32
timestamp 1490727624
transform 1 0 748 0 1 450
box -3 -3 3 3
use $$M2_M1  $$M2_M1_26
timestamp 1490727624
transform 1 0 740 0 1 440
box -2 -2 2 2
use $$M3_M2  $$M3_M2_33
timestamp 1490727624
transform 1 0 716 0 1 410
box -3 -3 3 3
use $$M3_M2  $$M3_M2_34
timestamp 1490727624
transform 1 0 740 0 1 410
box -3 -3 3 3
use $$M2_M1  $$M2_M1_27
timestamp 1490727624
transform 1 0 796 0 1 460
box -2 -2 2 2
use $$M3_M2  $$M3_M2_35
timestamp 1490727624
transform 1 0 796 0 1 450
box -3 -3 3 3
use $$M2_M1  $$M2_M1_28
timestamp 1490727624
transform 1 0 796 0 1 440
box -2 -2 2 2
use $$M3_M2  $$M3_M2_36
timestamp 1490727624
transform 1 0 796 0 1 440
box -3 -3 3 3
use $$M2_M1  $$M2_M1_29
timestamp 1490727624
transform 1 0 764 0 1 400
box -2 -2 2 2
use $$M2_M1  $$M2_M1_31
timestamp 1490727624
transform 1 0 900 0 1 450
box -2 -2 2 2
use $$M2_M1  $$M2_M1_30
timestamp 1490727624
transform 1 0 916 0 1 453
box -2 -2 2 2
use $$M3_M2  $$M3_M2_37
timestamp 1490727624
transform 1 0 900 0 1 440
box -3 -3 3 3
use $$M2_M1  $$M2_M1_32
timestamp 1490727624
transform 1 0 892 0 1 430
box -2 -2 2 2
use $$M3_M2  $$M3_M2_38
timestamp 1490727624
transform 1 0 924 0 1 400
box -3 -3 3 3
use $$M2_M1  $$M2_M1_33
timestamp 1490727624
transform 1 0 940 0 1 453
box -2 -2 2 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_1
timestamp 1490727624
transform 1 0 1009 0 1 490
box -7 -2 7 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_2
timestamp 1490727624
transform 1 0 37 0 1 390
box -7 -2 7 2
use FILL  FILL_0
timestamp 1490727624
transform 1 0 80 0 -1 490
box -8 -3 16 105
use NOR2X1  NOR2X1_0
timestamp 1490727624
transform -1 0 112 0 -1 490
box -8 -3 32 105
use FILL  FILL_1
timestamp 1490727624
transform 1 0 112 0 -1 490
box -8 -3 16 105
use OAI21X1  OAI21X1_0
timestamp 1490727624
transform 1 0 120 0 -1 490
box -8 -3 34 105
use FILL  FILL_2
timestamp 1490727624
transform 1 0 152 0 -1 490
box -8 -3 16 105
use FILL  FILL_3
timestamp 1490727624
transform 1 0 160 0 -1 490
box -8 -3 16 105
use $$M3_M2  $$M3_M2_39
timestamp 1490727624
transform 1 0 180 0 1 390
box -3 -3 3 3
use INVX2  INVX2_0
timestamp 1490727624
transform -1 0 184 0 -1 490
box -9 -3 26 105
use INVX2  INVX2_1
timestamp 1490727624
transform -1 0 200 0 -1 490
box -9 -3 26 105
use FILL  FILL_4
timestamp 1490727624
transform 1 0 200 0 -1 490
box -8 -3 16 105
use $$M3_M2  $$M3_M2_40
timestamp 1490727624
transform 1 0 220 0 1 390
box -3 -3 3 3
use FILL  FILL_5
timestamp 1490727624
transform 1 0 208 0 -1 490
box -8 -3 16 105
use DFFPOSX1  DFFPOSX1_0
timestamp 1490727624
transform -1 0 312 0 -1 490
box -8 -3 104 105
use FILL  FILL_6
timestamp 1490727624
transform 1 0 312 0 -1 490
box -8 -3 16 105
use FILL  FILL_7
timestamp 1490727624
transform 1 0 320 0 -1 490
box -8 -3 16 105
use FILL  FILL_8
timestamp 1490727624
transform 1 0 328 0 -1 490
box -8 -3 16 105
use FILL  FILL_9
timestamp 1490727624
transform 1 0 336 0 -1 490
box -8 -3 16 105
use FILL  FILL_10
timestamp 1490727624
transform 1 0 344 0 -1 490
box -8 -3 16 105
use FILL  FILL_11
timestamp 1490727624
transform 1 0 352 0 -1 490
box -8 -3 16 105
use FILL  FILL_12
timestamp 1490727624
transform 1 0 360 0 -1 490
box -8 -3 16 105
use FILL  FILL_13
timestamp 1490727624
transform 1 0 368 0 -1 490
box -8 -3 16 105
use DFFPOSX1  DFFPOSX1_1
timestamp 1490727624
transform -1 0 472 0 -1 490
box -8 -3 104 105
use FILL  FILL_14
timestamp 1490727624
transform 1 0 472 0 -1 490
box -8 -3 16 105
use FILL  FILL_15
timestamp 1490727624
transform 1 0 480 0 -1 490
box -8 -3 16 105
use AND2X2  AND2X2_0
timestamp 1490727624
transform 1 0 488 0 -1 490
box -8 -3 40 105
use FILL  FILL_16
timestamp 1490727624
transform 1 0 520 0 -1 490
box -8 -3 16 105
use INVX2  INVX2_2
timestamp 1490727624
transform -1 0 544 0 -1 490
box -9 -3 26 105
use FILL  FILL_17
timestamp 1490727624
transform 1 0 544 0 -1 490
box -8 -3 16 105
use FILL  FILL_18
timestamp 1490727624
transform 1 0 552 0 -1 490
box -8 -3 16 105
use DFFPOSX1  DFFPOSX1_2
timestamp 1490727624
transform -1 0 656 0 -1 490
box -8 -3 104 105
use FILL  FILL_19
timestamp 1490727624
transform 1 0 656 0 -1 490
box -8 -3 16 105
use FILL  FILL_20
timestamp 1490727624
transform 1 0 664 0 -1 490
box -8 -3 16 105
use AND2X2  AND2X2_1
timestamp 1490727624
transform -1 0 704 0 -1 490
box -8 -3 40 105
use LATCH  LATCH_0
timestamp 1490727624
transform -1 0 760 0 -1 490
box -8 -3 64 105
use LATCH  LATCH_1
timestamp 1490727624
transform -1 0 816 0 -1 490
box -8 -3 64 105
use FILL  FILL_21
timestamp 1490727624
transform 1 0 816 0 -1 490
box -8 -3 16 105
use FILL  FILL_22
timestamp 1490727624
transform 1 0 824 0 -1 490
box -8 -3 16 105
use FILL  FILL_23
timestamp 1490727624
transform 1 0 832 0 -1 490
box -8 -3 16 105
use FILL  FILL_24
timestamp 1490727624
transform 1 0 840 0 -1 490
box -8 -3 16 105
use FILL  FILL_25
timestamp 1490727624
transform 1 0 848 0 -1 490
box -8 -3 16 105
use FILL  FILL_26
timestamp 1490727624
transform 1 0 856 0 -1 490
box -8 -3 16 105
use FILL  FILL_27
timestamp 1490727624
transform 1 0 864 0 -1 490
box -8 -3 16 105
use FILL  FILL_28
timestamp 1490727624
transform 1 0 872 0 -1 490
box -8 -3 16 105
use FILL  FILL_29
timestamp 1490727624
transform 1 0 880 0 -1 490
box -8 -3 16 105
use OAI21X1  OAI21X1_1
timestamp 1490727624
transform -1 0 920 0 -1 490
box -8 -3 34 105
use FILL  FILL_30
timestamp 1490727624
transform 1 0 920 0 -1 490
box -8 -3 16 105
use INVX2  INVX2_3
timestamp 1490727624
transform -1 0 944 0 -1 490
box -9 -3 26 105
use FILL  FILL_31
timestamp 1490727624
transform 1 0 944 0 -1 490
box -8 -3 16 105
use FILL  FILL_32
timestamp 1490727624
transform 1 0 952 0 -1 490
box -8 -3 16 105
use FILL  FILL_33
timestamp 1490727624
transform 1 0 960 0 -1 490
box -8 -3 16 105
use FILL  FILL_34
timestamp 1490727624
transform 1 0 968 0 -1 490
box -8 -3 16 105
use FILL  FILL_35
timestamp 1490727624
transform 1 0 976 0 -1 490
box -8 -3 16 105
use FILL  FILL_36
timestamp 1490727624
transform 1 0 984 0 -1 490
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_3
timestamp 1490727624
transform 1 0 1034 0 1 390
box -7 -2 7 2
use $$M2_M1  $$M2_M1_34
timestamp 1490727624
transform 1 0 92 0 1 380
box -2 -2 2 2
use $$M2_M1  $$M2_M1_36
timestamp 1490727624
transform 1 0 100 0 1 350
box -2 -2 2 2
use $$M3_M2  $$M3_M2_41
timestamp 1490727624
transform 1 0 100 0 1 350
box -3 -3 3 3
use $$M2_M1  $$M2_M1_38
timestamp 1490727624
transform 1 0 84 0 1 321
box -2 -2 2 2
use $$M3_M2  $$M3_M2_43
timestamp 1490727624
transform 1 0 92 0 1 320
box -3 -3 3 3
use $$M2_M1  $$M2_M1_37
timestamp 1490727624
transform 1 0 116 0 1 350
box -2 -2 2 2
use $$M3_M2  $$M3_M2_42
timestamp 1490727624
transform 1 0 116 0 1 330
box -3 -3 3 3
use $$M2_M1  $$M2_M1_35
timestamp 1490727624
transform 1 0 132 0 1 380
box -2 -2 2 2
use $$M2_M1  $$M2_M1_39
timestamp 1490727624
transform 1 0 161 0 1 360
box -2 -2 2 2
use $$M3_M2  $$M3_M2_44
timestamp 1490727624
transform 1 0 161 0 1 360
box -3 -3 3 3
use $$M2_M1  $$M2_M1_42
timestamp 1490727624
transform 1 0 164 0 1 339
box -2 -2 2 2
use $$M3_M2  $$M3_M2_47
timestamp 1490727624
transform 1 0 156 0 1 330
box -3 -3 3 3
use $$M2_M1  $$M2_M1_44
timestamp 1490727624
transform 1 0 148 0 1 323
box -2 -2 2 2
use $$M2_M1  $$M2_M1_45
timestamp 1490727624
transform 1 0 148 0 1 315
box -2 -2 2 2
use $$M2_M1  $$M2_M1_46
timestamp 1490727624
transform 1 0 180 0 1 320
box -2 -2 2 2
use $$M3_M2  $$M3_M2_49
timestamp 1490727624
transform 1 0 180 0 1 320
box -3 -3 3 3
use $$M3_M2  $$M3_M2_45
timestamp 1490727624
transform 1 0 204 0 1 360
box -3 -3 3 3
use $$M2_M1  $$M2_M1_40
timestamp 1490727624
transform 1 0 196 0 1 350
box -2 -2 2 2
use $$M2_M1  $$M2_M1_41
timestamp 1490727624
transform 1 0 204 0 1 350
box -2 -2 2 2
use $$M3_M2  $$M3_M2_46
timestamp 1490727624
transform 1 0 204 0 1 340
box -3 -3 3 3
use $$M2_M1  $$M2_M1_43
timestamp 1490727624
transform 1 0 204 0 1 335
box -2 -2 2 2
use $$M3_M2  $$M3_M2_48
timestamp 1490727624
transform 1 0 212 0 1 330
box -3 -3 3 3
use $$M3_M2  $$M3_M2_50
timestamp 1490727624
transform 1 0 228 0 1 360
box -3 -3 3 3
use $$M2_M1  $$M2_M1_47
timestamp 1490727624
transform 1 0 228 0 1 327
box -2 -2 2 2
use $$M3_M2  $$M3_M2_51
timestamp 1490727624
transform 1 0 244 0 1 340
box -3 -3 3 3
use $$M2_M1  $$M2_M1_48
timestamp 1490727624
transform 1 0 244 0 1 327
box -2 -2 2 2
use $$M2_M1  $$M2_M1_49
timestamp 1490727624
transform 1 0 236 0 1 310
box -2 -2 2 2
use $$M3_M2  $$M3_M2_52
timestamp 1490727624
transform 1 0 236 0 1 310
box -3 -3 3 3
use $$M2_M1  $$M2_M1_51
timestamp 1490727624
transform 1 0 276 0 1 380
box -2 -2 2 2
use $$M2_M1  $$M2_M1_57
timestamp 1490727624
transform 1 0 268 0 1 311
box -2 -2 2 2
use $$M3_M2  $$M3_M2_56
timestamp 1490727624
transform 1 0 268 0 1 310
box -3 -3 3 3
use $$M2_M1  $$M2_M1_50
timestamp 1490727624
transform 1 0 252 0 1 300
box -2 -2 2 2
use $$M3_M2  $$M3_M2_53
timestamp 1490727624
transform 1 0 300 0 1 380
box -3 -3 3 3
use $$M2_M1  $$M2_M1_54
timestamp 1490727624
transform 1 0 292 0 1 333
box -2 -2 2 2
use $$M2_M1  $$M2_M1_52
timestamp 1490727624
transform 1 0 322 0 1 380
box -2 -2 2 2
use $$M3_M2  $$M3_M2_55
timestamp 1490727624
transform 1 0 308 0 1 340
box -3 -3 3 3
use $$M3_M2  $$M3_M2_54
timestamp 1490727624
transform 1 0 332 0 1 350
box -3 -3 3 3
use $$M2_M1  $$M2_M1_53
timestamp 1490727624
transform 1 0 332 0 1 344
box -2 -2 2 2
use $$M2_M1  $$M2_M1_55
timestamp 1490727624
transform 1 0 316 0 1 331
box -2 -2 2 2
use $$M2_M1  $$M2_M1_56
timestamp 1490727624
transform 1 0 308 0 1 327
box -2 -2 2 2
use $$M3_M2  $$M3_M2_58
timestamp 1490727624
transform 1 0 300 0 1 300
box -3 -3 3 3
use $$M3_M2  $$M3_M2_57
timestamp 1490727624
transform 1 0 316 0 1 310
box -3 -3 3 3
use $$M3_M2  $$M3_M2_60
timestamp 1490727624
transform 1 0 348 0 1 330
box -3 -3 3 3
use $$M2_M1  $$M2_M1_59
timestamp 1490727624
transform 1 0 348 0 1 321
box -2 -2 2 2
use $$M2_M1  $$M2_M1_58
timestamp 1490727624
transform 1 0 364 0 1 380
box -2 -2 2 2
use $$M3_M2  $$M3_M2_59
timestamp 1490727624
transform 1 0 364 0 1 380
box -3 -3 3 3
use $$M3_M2  $$M3_M2_61
timestamp 1490727624
transform 1 0 356 0 1 310
box -3 -3 3 3
use $$M2_M1  $$M2_M1_60
timestamp 1490727624
transform 1 0 356 0 1 300
box -2 -2 2 2
use $$M3_M2  $$M3_M2_62
timestamp 1490727624
transform 1 0 380 0 1 340
box -3 -3 3 3
use $$M3_M2  $$M3_M2_64
timestamp 1490727624
transform 1 0 372 0 1 310
box -3 -3 3 3
use $$M2_M1  $$M2_M1_61
timestamp 1490727624
transform 1 0 396 0 1 330
box -2 -2 2 2
use $$M3_M2  $$M3_M2_63
timestamp 1490727624
transform 1 0 396 0 1 330
box -3 -3 3 3
use $$M2_M1  $$M2_M1_62
timestamp 1490727624
transform 1 0 404 0 1 330
box -2 -2 2 2
use $$M3_M2  $$M3_M2_67
timestamp 1490727624
transform 1 0 444 0 1 350
box -3 -3 3 3
use $$M3_M2  $$M3_M2_68
timestamp 1490727624
transform 1 0 428 0 1 340
box -3 -3 3 3
use $$M2_M1  $$M2_M1_63
timestamp 1490727624
transform 1 0 444 0 1 340
box -2 -2 2 2
use $$M3_M2  $$M3_M2_74
timestamp 1490727624
transform 1 0 420 0 1 320
box -3 -3 3 3
use $$M2_M1  $$M2_M1_68
timestamp 1490727624
transform 1 0 428 0 1 320
box -2 -2 2 2
use $$M2_M1  $$M2_M1_70
timestamp 1490727624
transform 1 0 420 0 1 312
box -2 -2 2 2
use $$M3_M2  $$M3_M2_75
timestamp 1490727624
transform 1 0 460 0 1 320
box -3 -3 3 3
use $$M2_M1  $$M2_M1_71
timestamp 1490727624
transform 1 0 460 0 1 310
box -2 -2 2 2
use $$M3_M2  $$M3_M2_66
timestamp 1490727624
transform 1 0 548 0 1 360
box -3 -3 3 3
use $$M2_M1  $$M2_M1_69
timestamp 1490727624
transform 1 0 532 0 1 320
box -2 -2 2 2
use $$M3_M2  $$M3_M2_69
timestamp 1490727624
transform 1 0 564 0 1 340
box -3 -3 3 3
use $$M3_M2  $$M3_M2_76
timestamp 1490727624
transform 1 0 564 0 1 320
box -3 -3 3 3
use $$M3_M2  $$M3_M2_65
timestamp 1490727624
transform 1 0 604 0 1 370
box -3 -3 3 3
use $$M2_M1  $$M2_M1_65
timestamp 1490727624
transform 1 0 596 0 1 330
box -2 -2 2 2
use $$M3_M2  $$M3_M2_72
timestamp 1490727624
transform 1 0 596 0 1 330
box -3 -3 3 3
use $$M3_M2  $$M3_M2_70
timestamp 1490727624
transform 1 0 612 0 1 340
box -3 -3 3 3
use $$M2_M1  $$M2_M1_66
timestamp 1490727624
transform 1 0 604 0 1 330
box -2 -2 2 2
use $$M3_M2  $$M3_M2_71
timestamp 1490727624
transform 1 0 644 0 1 340
box -3 -3 3 3
use $$M2_M1  $$M2_M1_67
timestamp 1490727624
transform 1 0 636 0 1 330
box -2 -2 2 2
use $$M3_M2  $$M3_M2_73
timestamp 1490727624
transform 1 0 636 0 1 330
box -3 -3 3 3
use $$M2_M1  $$M2_M1_64
timestamp 1490727624
transform 1 0 644 0 1 333
box -2 -2 2 2
use $$M2_M1  $$M2_M1_75
timestamp 1490727624
transform 1 0 628 0 1 319
box -2 -2 2 2
use $$M3_M2  $$M3_M2_79
timestamp 1490727624
transform 1 0 628 0 1 320
box -3 -3 3 3
use $$M2_M1  $$M2_M1_74
timestamp 1490727624
transform 1 0 652 0 1 323
box -2 -2 2 2
use $$M3_M2  $$M3_M2_77
timestamp 1490727624
transform 1 0 668 0 1 340
box -3 -3 3 3
use $$M2_M1  $$M2_M1_72
timestamp 1490727624
transform 1 0 681 0 1 344
box -2 -2 2 2
use $$M2_M1  $$M2_M1_73
timestamp 1490727624
transform 1 0 668 0 1 331
box -2 -2 2 2
use $$M3_M2  $$M3_M2_78
timestamp 1490727624
transform 1 0 681 0 1 330
box -3 -3 3 3
use $$M2_M1  $$M2_M1_76
timestamp 1490727624
transform 1 0 716 0 1 380
box -2 -2 2 2
use $$M2_M1  $$M2_M1_78
timestamp 1490727624
transform 1 0 732 0 1 340
box -2 -2 2 2
use $$M3_M2  $$M3_M2_81
timestamp 1490727624
transform 1 0 732 0 1 340
box -3 -3 3 3
use $$M3_M2  $$M3_M2_80
timestamp 1490727624
transform 1 0 764 0 1 370
box -3 -3 3 3
use $$M3_M2  $$M3_M2_82
timestamp 1490727624
transform 1 0 756 0 1 330
box -3 -3 3 3
use $$M2_M1  $$M2_M1_81
timestamp 1490727624
transform 1 0 748 0 1 320
box -2 -2 2 2
use $$M2_M1  $$M2_M1_82
timestamp 1490727624
transform 1 0 756 0 1 317
box -2 -2 2 2
use $$M2_M1  $$M2_M1_77
timestamp 1490727624
transform 1 0 796 0 1 350
box -2 -2 2 2
use $$M2_M1  $$M2_M1_79
timestamp 1490727624
transform 1 0 788 0 1 340
box -2 -2 2 2
use $$M3_M2  $$M3_M2_83
timestamp 1490727624
transform 1 0 788 0 1 330
box -3 -3 3 3
use $$M2_M1  $$M2_M1_80
timestamp 1490727624
transform 1 0 780 0 1 322
box -2 -2 2 2
use $$M3_M2  $$M3_M2_84
timestamp 1490727624
transform 1 0 780 0 1 320
box -3 -3 3 3
use $$M3_M2  $$M3_M2_86
timestamp 1490727624
transform 1 0 820 0 1 360
box -3 -3 3 3
use $$M2_M1  $$M2_M1_85
timestamp 1490727624
transform 1 0 828 0 1 350
box -2 -2 2 2
use $$M2_M1  $$M2_M1_86
timestamp 1490727624
transform 1 0 812 0 1 340
box -2 -2 2 2
use $$M3_M2  $$M3_M2_88
timestamp 1490727624
transform 1 0 812 0 1 330
box -3 -3 3 3
use $$M2_M1  $$M2_M1_87
timestamp 1490727624
transform 1 0 820 0 1 334
box -2 -2 2 2
use $$M2_M1  $$M2_M1_89
timestamp 1490727624
transform 1 0 836 0 1 330
box -2 -2 2 2
use $$M3_M2  $$M3_M2_89
timestamp 1490727624
transform 1 0 836 0 1 330
box -3 -3 3 3
use $$M3_M2  $$M3_M2_91
timestamp 1490727624
transform 1 0 828 0 1 300
box -3 -3 3 3
use $$M2_M1  $$M2_M1_84
timestamp 1490727624
transform 1 0 863 0 1 370
box -2 -2 2 2
use $$M3_M2  $$M3_M2_85
timestamp 1490727624
transform 1 0 863 0 1 370
box -3 -3 3 3
use $$M2_M1  $$M2_M1_88
timestamp 1490727624
transform 1 0 860 0 1 333
box -2 -2 2 2
use $$M3_M2  $$M3_M2_90
timestamp 1490727624
transform 1 0 860 0 1 320
box -3 -3 3 3
use $$M3_M2  $$M3_M2_87
timestamp 1490727624
transform 1 0 876 0 1 350
box -3 -3 3 3
use $$M2_M1  $$M2_M1_90
timestamp 1490727624
transform 1 0 876 0 1 311
box -2 -2 2 2
use $$M2_M1  $$M2_M1_83
timestamp 1490727624
transform 1 0 892 0 1 380
box -2 -2 2 2
use $$M3_M2  $$M3_M2_92
timestamp 1490727624
transform 1 0 940 0 1 370
box -3 -3 3 3
use $$M2_M1  $$M2_M1_91
timestamp 1490727624
transform 1 0 948 0 1 330
box -2 -2 2 2
use $$M3_M2  $$M3_M2_93
timestamp 1490727624
transform 1 0 948 0 1 330
box -3 -3 3 3
use $$M2_M1  $$M2_M1_92
timestamp 1490727624
transform 1 0 956 0 1 330
box -2 -2 2 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_4
timestamp 1490727624
transform 1 0 62 0 1 290
box -7 -2 7 2
use NAND2X1  NAND2X1_0
timestamp 1490727624
transform 1 0 80 0 1 290
box -8 -3 32 105
use FILL  FILL_37
timestamp 1490727624
transform -1 0 112 0 1 290
box -8 -3 16 105
use FILL  FILL_38
timestamp 1490727624
transform -1 0 120 0 1 290
box -8 -3 16 105
use NAND2X1  NAND2X1_1
timestamp 1490727624
transform -1 0 144 0 1 290
box -8 -3 32 105
use $$M3_M2  $$M3_M2_94
timestamp 1490727624
transform 1 0 172 0 1 290
box -3 -3 3 3
use NOR2X1  NOR2X1_1
timestamp 1490727624
transform 1 0 144 0 1 290
box -8 -3 32 105
use FILL  FILL_42
timestamp 1490727624
transform -1 0 176 0 1 290
box -8 -3 16 105
use FILL  FILL_43
timestamp 1490727624
transform -1 0 184 0 1 290
box -8 -3 16 105
use NAND3X1  NAND3X1_0
timestamp 1490727624
transform -1 0 216 0 1 290
box -8 -3 40 105
use FILL  FILL_47
timestamp 1490727624
transform -1 0 224 0 1 290
box -8 -3 16 105
use INVX2  INVX2_4
timestamp 1490727624
transform 1 0 224 0 1 290
box -9 -3 26 105
use INVX2  INVX2_5
timestamp 1490727624
transform 1 0 240 0 1 290
box -9 -3 26 105
use FILL  FILL_49
timestamp 1490727624
transform -1 0 264 0 1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_2
timestamp 1490727624
transform 1 0 264 0 1 290
box -8 -3 32 105
use FILL  FILL_50
timestamp 1490727624
transform -1 0 296 0 1 290
box -8 -3 16 105
use FILL  FILL_51
timestamp 1490727624
transform -1 0 304 0 1 290
box -8 -3 16 105
use OAI21X1  OAI21X1_2
timestamp 1490727624
transform 1 0 304 0 1 290
box -8 -3 34 105
use FILL  FILL_54
timestamp 1490727624
transform -1 0 344 0 1 290
box -8 -3 16 105
use INVX2  INVX2_6
timestamp 1490727624
transform 1 0 344 0 1 290
box -9 -3 26 105
use FILL  FILL_56
timestamp 1490727624
transform -1 0 368 0 1 290
box -8 -3 16 105
use FILL  FILL_58
timestamp 1490727624
transform -1 0 376 0 1 290
box -8 -3 16 105
use AND2X2  AND2X2_2
timestamp 1490727624
transform -1 0 408 0 1 290
box -8 -3 40 105
use FILL  FILL_59
timestamp 1490727624
transform -1 0 416 0 1 290
box -8 -3 16 105
use OR2X1  OR2X1_0
timestamp 1490727624
transform 1 0 416 0 1 290
box -8 -3 40 105
use FILL  FILL_60
timestamp 1490727624
transform -1 0 456 0 1 290
box -8 -3 16 105
use FILL  FILL_61
timestamp 1490727624
transform -1 0 464 0 1 290
box -8 -3 16 105
use DFFPOSX1  DFFPOSX1_3
timestamp 1490727624
transform -1 0 560 0 1 290
box -8 -3 104 105
use FILL  FILL_62
timestamp 1490727624
transform -1 0 568 0 1 290
box -8 -3 16 105
use FILL  FILL_63
timestamp 1490727624
transform -1 0 576 0 1 290
box -8 -3 16 105
use AND2X2  AND2X2_3
timestamp 1490727624
transform -1 0 608 0 1 290
box -8 -3 40 105
use FILL  FILL_64
timestamp 1490727624
transform -1 0 616 0 1 290
box -8 -3 16 105
use FILL  FILL_65
timestamp 1490727624
transform -1 0 624 0 1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_3
timestamp 1490727624
transform 1 0 624 0 1 290
box -8 -3 32 105
use FILL  FILL_74
timestamp 1490727624
transform -1 0 656 0 1 290
box -8 -3 16 105
use OAI21X1  OAI21X1_3
timestamp 1490727624
transform 1 0 656 0 1 290
box -8 -3 34 105
use FILL  FILL_76
timestamp 1490727624
transform -1 0 696 0 1 290
box -8 -3 16 105
use FILL  FILL_77
timestamp 1490727624
transform -1 0 704 0 1 290
box -8 -3 16 105
use INVX2  INVX2_7
timestamp 1490727624
transform 1 0 704 0 1 290
box -9 -3 26 105
use FILL  FILL_79
timestamp 1490727624
transform -1 0 728 0 1 290
box -8 -3 16 105
use OR2X1  OR2X1_1
timestamp 1490727624
transform -1 0 760 0 1 290
box -8 -3 40 105
use FILL  FILL_81
timestamp 1490727624
transform -1 0 768 0 1 290
box -8 -3 16 105
use FILL  FILL_82
timestamp 1490727624
transform -1 0 776 0 1 290
box -8 -3 16 105
use NAND2X1  NAND2X1_2
timestamp 1490727624
transform 1 0 776 0 1 290
box -8 -3 32 105
use FILL  FILL_83
timestamp 1490727624
transform -1 0 808 0 1 290
box -8 -3 16 105
use NAND3X1  NAND3X1_1
timestamp 1490727624
transform 1 0 808 0 1 290
box -8 -3 40 105
use FILL  FILL_84
timestamp 1490727624
transform -1 0 848 0 1 290
box -8 -3 16 105
use FILL  FILL_85
timestamp 1490727624
transform -1 0 856 0 1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_4
timestamp 1490727624
transform -1 0 880 0 1 290
box -8 -3 32 105
use FILL  FILL_93
timestamp 1490727624
transform -1 0 888 0 1 290
box -8 -3 16 105
use FILL  FILL_94
timestamp 1490727624
transform -1 0 896 0 1 290
box -8 -3 16 105
use FILL  FILL_95
timestamp 1490727624
transform -1 0 904 0 1 290
box -8 -3 16 105
use FILL  FILL_96
timestamp 1490727624
transform -1 0 912 0 1 290
box -8 -3 16 105
use FILL  FILL_97
timestamp 1490727624
transform -1 0 920 0 1 290
box -8 -3 16 105
use FILL  FILL_98
timestamp 1490727624
transform -1 0 928 0 1 290
box -8 -3 16 105
use AND2X2  AND2X2_4
timestamp 1490727624
transform -1 0 960 0 1 290
box -8 -3 40 105
use FILL  FILL_101
timestamp 1490727624
transform -1 0 968 0 1 290
box -8 -3 16 105
use FILL  FILL_102
timestamp 1490727624
transform -1 0 976 0 1 290
box -8 -3 16 105
use FILL  FILL_103
timestamp 1490727624
transform -1 0 984 0 1 290
box -8 -3 16 105
use FILL  FILL_104
timestamp 1490727624
transform -1 0 992 0 1 290
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_6
timestamp 1490727624
transform 1 0 1009 0 1 290
box -7 -2 7 2
use $$M2_M1  $$M2_M1_93
timestamp 1490727624
transform 1 0 92 0 1 259
box -2 -2 2 2
use $$M3_M2  $$M3_M2_95
timestamp 1490727624
transform 1 0 20 0 1 200
box -3 -3 3 3
use $$M2_M1  $$M2_M1_94
timestamp 1490727624
transform 1 0 84 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_96
timestamp 1490727624
transform 1 0 84 0 1 200
box -3 -3 3 3
use $$M3_M2  $$M3_M2_97
timestamp 1490727624
transform 1 0 108 0 1 280
box -3 -3 3 3
use $$M3_M2  $$M3_M2_98
timestamp 1490727624
transform 1 0 108 0 1 210
box -3 -3 3 3
use $$M2_M1  $$M2_M1_95
timestamp 1490727624
transform 1 0 108 0 1 200
box -2 -2 2 2
use $$M2_M1  $$M2_M1_98
timestamp 1490727624
transform 1 0 156 0 1 244
box -2 -2 2 2
use $$M3_M2  $$M3_M2_102
timestamp 1490727624
transform 1 0 156 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_99
timestamp 1490727624
transform 1 0 164 0 1 240
box -2 -2 2 2
use $$M2_M1  $$M2_M1_101
timestamp 1490727624
transform 1 0 148 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_104
timestamp 1490727624
transform 1 0 148 0 1 230
box -3 -3 3 3
use $$M3_M2  $$M3_M2_105
timestamp 1490727624
transform 1 0 164 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_106
timestamp 1490727624
transform 1 0 172 0 1 210
box -3 -3 3 3
use $$M2_M1  $$M2_M1_96
timestamp 1490727624
transform 1 0 196 0 1 270
box -2 -2 2 2
use $$M3_M2  $$M3_M2_99
timestamp 1490727624
transform 1 0 196 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_97
timestamp 1490727624
transform 1 0 188 0 1 264
box -2 -2 2 2
use $$M3_M2  $$M3_M2_100
timestamp 1490727624
transform 1 0 188 0 1 260
box -3 -3 3 3
use $$M3_M2  $$M3_M2_107
timestamp 1490727624
transform 1 0 188 0 1 210
box -3 -3 3 3
use $$M3_M2  $$M3_M2_101
timestamp 1490727624
transform 1 0 204 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_100
timestamp 1490727624
transform 1 0 204 0 1 241
box -2 -2 2 2
use $$M3_M2  $$M3_M2_103
timestamp 1490727624
transform 1 0 204 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_102
timestamp 1490727624
transform 1 0 220 0 1 280
box -2 -2 2 2
use $$M3_M2  $$M3_M2_108
timestamp 1490727624
transform 1 0 244 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_103
timestamp 1490727624
transform 1 0 244 0 1 256
box -2 -2 2 2
use $$M3_M2  $$M3_M2_109
timestamp 1490727624
transform 1 0 236 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_104
timestamp 1490727624
transform 1 0 244 0 1 242
box -2 -2 2 2
use $$M2_M1  $$M2_M1_105
timestamp 1490727624
transform 1 0 222 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_110
timestamp 1490727624
transform 1 0 222 0 1 230
box -3 -3 3 3
use $$M3_M2  $$M3_M2_111
timestamp 1490727624
transform 1 0 244 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_112
timestamp 1490727624
transform 1 0 268 0 1 280
box -3 -3 3 3
use $$M3_M2  $$M3_M2_113
timestamp 1490727624
transform 1 0 268 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_109
timestamp 1490727624
transform 1 0 260 0 1 230
box -2 -2 2 2
use $$M2_M1  $$M2_M1_107
timestamp 1490727624
transform 1 0 284 0 1 260
box -2 -2 2 2
use $$M2_M1  $$M2_M1_108
timestamp 1490727624
transform 1 0 276 0 1 253
box -2 -2 2 2
use $$M3_M2  $$M3_M2_114
timestamp 1490727624
transform 1 0 276 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_110
timestamp 1490727624
transform 1 0 268 0 1 200
box -2 -2 2 2
use $$M2_M1  $$M2_M1_106
timestamp 1490727624
transform 1 0 300 0 1 280
box -2 -2 2 2
use $$M3_M2  $$M3_M2_115
timestamp 1490727624
transform 1 0 292 0 1 220
box -3 -3 3 3
use $$M2_M1  $$M2_M1_111
timestamp 1490727624
transform 1 0 332 0 1 263
box -2 -2 2 2
use $$M3_M2  $$M3_M2_116
timestamp 1490727624
transform 1 0 332 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_112
timestamp 1490727624
transform 1 0 316 0 1 241
box -2 -2 2 2
use $$M2_M1  $$M2_M1_113
timestamp 1490727624
transform 1 0 324 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_117
timestamp 1490727624
transform 1 0 324 0 1 240
box -3 -3 3 3
use $$M3_M2  $$M3_M2_118
timestamp 1490727624
transform 1 0 316 0 1 220
box -3 -3 3 3
use $$M2_M1  $$M2_M1_114
timestamp 1490727624
transform 1 0 356 0 1 263
box -2 -2 2 2
use $$M3_M2  $$M3_M2_119
timestamp 1490727624
transform 1 0 356 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_115
timestamp 1490727624
transform 1 0 348 0 1 200
box -2 -2 2 2
use $$M2_M1  $$M2_M1_116
timestamp 1490727624
transform 1 0 380 0 1 260
box -2 -2 2 2
use $$M3_M2  $$M3_M2_120
timestamp 1490727624
transform 1 0 380 0 1 260
box -3 -3 3 3
use $$M3_M2  $$M3_M2_121
timestamp 1490727624
transform 1 0 404 0 1 280
box -3 -3 3 3
use $$M2_M1  $$M2_M1_117
timestamp 1490727624
transform 1 0 444 0 1 280
box -2 -2 2 2
use $$M3_M2  $$M3_M2_122
timestamp 1490727624
transform 1 0 444 0 1 280
box -3 -3 3 3
use $$M2_M1  $$M2_M1_119
timestamp 1490727624
transform 1 0 388 0 1 259
box -2 -2 2 2
use $$M2_M1  $$M2_M1_118
timestamp 1490727624
transform 1 0 412 0 1 260
box -2 -2 2 2
use $$M2_M1  $$M2_M1_121
timestamp 1490727624
transform 1 0 372 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_123
timestamp 1490727624
transform 1 0 412 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_120
timestamp 1490727624
transform 1 0 412 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_124
timestamp 1490727624
transform 1 0 388 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_122
timestamp 1490727624
transform 1 0 380 0 1 200
box -2 -2 2 2
use $$M2_M1  $$M2_M1_123
timestamp 1490727624
transform 1 0 460 0 1 280
box -2 -2 2 2
use $$M3_M2  $$M3_M2_125
timestamp 1490727624
transform 1 0 460 0 1 280
box -3 -3 3 3
use $$M3_M2  $$M3_M2_126
timestamp 1490727624
transform 1 0 484 0 1 280
box -3 -3 3 3
use $$M2_M1  $$M2_M1_124
timestamp 1490727624
transform 1 0 500 0 1 255
box -2 -2 2 2
use $$M3_M2  $$M3_M2_127
timestamp 1490727624
transform 1 0 500 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_125
timestamp 1490727624
transform 1 0 492 0 1 230
box -2 -2 2 2
use $$M2_M1  $$M2_M1_126
timestamp 1490727624
transform 1 0 516 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_128
timestamp 1490727624
transform 1 0 572 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_127
timestamp 1490727624
transform 1 0 556 0 1 263
box -2 -2 2 2
use $$M2_M1  $$M2_M1_128
timestamp 1490727624
transform 1 0 572 0 1 251
box -2 -2 2 2
use $$M3_M2  $$M3_M2_129
timestamp 1490727624
transform 1 0 556 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_129
timestamp 1490727624
transform 1 0 580 0 1 243
box -2 -2 2 2
use $$M3_M2  $$M3_M2_131
timestamp 1490727624
transform 1 0 596 0 1 220
box -3 -3 3 3
use $$M2_M1  $$M2_M1_130
timestamp 1490727624
transform 1 0 612 0 1 263
box -2 -2 2 2
use $$M3_M2  $$M3_M2_130
timestamp 1490727624
transform 1 0 612 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_131
timestamp 1490727624
transform 1 0 628 0 1 241
box -2 -2 2 2
use $$M3_M2  $$M3_M2_132
timestamp 1490727624
transform 1 0 628 0 1 220
box -3 -3 3 3
use $$M2_M1  $$M2_M1_132
timestamp 1490727624
transform 1 0 625 0 1 210
box -2 -2 2 2
use $$M3_M2  $$M3_M2_133
timestamp 1490727624
transform 1 0 625 0 1 210
box -3 -3 3 3
use $$M3_M2  $$M3_M2_134
timestamp 1490727624
transform 1 0 652 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_135
timestamp 1490727624
transform 1 0 660 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_135
timestamp 1490727624
transform 1 0 652 0 1 230
box -2 -2 2 2
use $$M2_M1  $$M2_M1_136
timestamp 1490727624
transform 1 0 660 0 1 200
box -2 -2 2 2
use $$M2_M1  $$M2_M1_134
timestamp 1490727624
transform 1 0 676 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_136
timestamp 1490727624
transform 1 0 708 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_133
timestamp 1490727624
transform 1 0 700 0 1 243
box -2 -2 2 2
use $$M2_M1  $$M2_M1_137
timestamp 1490727624
transform 1 0 692 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_137
timestamp 1490727624
transform 1 0 692 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_138
timestamp 1490727624
transform 1 0 740 0 1 253
box -2 -2 2 2
use $$M3_M2  $$M3_M2_138
timestamp 1490727624
transform 1 0 740 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_139
timestamp 1490727624
transform 1 0 748 0 1 250
box -2 -2 2 2
use $$M3_M2  $$M3_M2_139
timestamp 1490727624
transform 1 0 740 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_140
timestamp 1490727624
transform 1 0 788 0 1 280
box -2 -2 2 2
use $$M2_M1  $$M2_M1_141
timestamp 1490727624
transform 1 0 804 0 1 255
box -2 -2 2 2
use $$M2_M1  $$M2_M1_143
timestamp 1490727624
transform 1 0 796 0 1 200
box -2 -2 2 2
use $$M2_M1  $$M2_M1_142
timestamp 1490727624
transform 1 0 812 0 1 250
box -2 -2 2 2
use $$M3_M2  $$M3_M2_140
timestamp 1490727624
transform 1 0 820 0 1 280
box -3 -3 3 3
use $$M2_M1  $$M2_M1_148
timestamp 1490727624
transform 1 0 836 0 1 249
box -2 -2 2 2
use $$M3_M2  $$M3_M2_141
timestamp 1490727624
transform 1 0 884 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_146
timestamp 1490727624
transform 1 0 860 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_147
timestamp 1490727624
transform 1 0 868 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_149
timestamp 1490727624
transform 1 0 852 0 1 233
box -2 -2 2 2
use $$M3_M2  $$M3_M2_145
timestamp 1490727624
transform 1 0 852 0 1 210
box -3 -3 3 3
use $$M3_M2  $$M3_M2_144
timestamp 1490727624
transform 1 0 876 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_150
timestamp 1490727624
transform 1 0 884 0 1 249
box -2 -2 2 2
use $$M3_M2  $$M3_M2_146
timestamp 1490727624
transform 1 0 868 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_151
timestamp 1490727624
transform 1 0 868 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_142
timestamp 1490727624
transform 1 0 916 0 1 280
box -3 -3 3 3
use $$M3_M2  $$M3_M2_143
timestamp 1490727624
transform 1 0 924 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_145
timestamp 1490727624
transform 1 0 900 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_144
timestamp 1490727624
transform 1 0 908 0 1 256
box -2 -2 2 2
use $$M3_M2  $$M3_M2_148
timestamp 1490727624
transform 1 0 900 0 1 210
box -3 -3 3 3
use $$M2_M1  $$M2_M1_152
timestamp 1490727624
transform 1 0 916 0 1 243
box -2 -2 2 2
use $$M3_M2  $$M3_M2_147
timestamp 1490727624
transform 1 0 916 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_153
timestamp 1490727624
transform 1 0 932 0 1 230
box -2 -2 2 2
use $$M2_M1  $$M2_M1_154
timestamp 1490727624
transform 1 0 948 0 1 280
box -2 -2 2 2
use $$M3_M2  $$M3_M2_151
timestamp 1490727624
transform 1 0 956 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_156
timestamp 1490727624
transform 1 0 956 0 1 247
box -2 -2 2 2
use $$M3_M2  $$M3_M2_149
timestamp 1490727624
transform 1 0 972 0 1 280
box -3 -3 3 3
use $$M2_M1  $$M2_M1_155
timestamp 1490727624
transform 1 0 972 0 1 260
box -2 -2 2 2
use $$M3_M2  $$M3_M2_150
timestamp 1490727624
transform 1 0 972 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_157
timestamp 1490727624
transform 1 0 959 0 1 200
box -2 -2 2 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_5
timestamp 1490727624
transform 1 0 37 0 1 190
box -7 -2 7 2
use INVX2  INVX2_8
timestamp 1490727624
transform -1 0 96 0 -1 290
box -9 -3 26 105
use FILL  FILL_39
timestamp 1490727624
transform 1 0 96 0 -1 290
box -8 -3 16 105
use INVX2  INVX2_9
timestamp 1490727624
transform -1 0 120 0 -1 290
box -9 -3 26 105
use FILL  FILL_40
timestamp 1490727624
transform 1 0 120 0 -1 290
box -8 -3 16 105
use FILL  FILL_41
timestamp 1490727624
transform 1 0 128 0 -1 290
box -8 -3 16 105
use NAND3X1  NAND3X1_2
timestamp 1490727624
transform -1 0 168 0 -1 290
box -8 -3 40 105
use FILL  FILL_44
timestamp 1490727624
transform 1 0 168 0 -1 290
box -8 -3 16 105
use FILL  FILL_45
timestamp 1490727624
transform 1 0 176 0 -1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_5
timestamp 1490727624
transform 1 0 184 0 -1 290
box -8 -3 32 105
use FILL  FILL_46
timestamp 1490727624
transform 1 0 208 0 -1 290
box -8 -3 16 105
use OAI21X1  OAI21X1_4
timestamp 1490727624
transform -1 0 248 0 -1 290
box -8 -3 34 105
use FILL  FILL_48
timestamp 1490727624
transform 1 0 248 0 -1 290
box -8 -3 16 105
use NAND2X1  NAND2X1_3
timestamp 1490727624
transform -1 0 280 0 -1 290
box -8 -3 32 105
use FILL  FILL_52
timestamp 1490727624
transform 1 0 280 0 -1 290
box -8 -3 16 105
use $$M3_M2  $$M3_M2_152
timestamp 1490727624
transform 1 0 316 0 1 190
box -3 -3 3 3
use INVX2  INVX2_10
timestamp 1490727624
transform 1 0 288 0 -1 290
box -9 -3 26 105
use FILL  FILL_53
timestamp 1490727624
transform 1 0 304 0 -1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_6
timestamp 1490727624
transform -1 0 336 0 -1 290
box -8 -3 32 105
use FILL  FILL_55
timestamp 1490727624
transform 1 0 336 0 -1 290
box -8 -3 16 105
use INVX1  INVX1_0
timestamp 1490727624
transform -1 0 360 0 -1 290
box -9 -3 26 105
use FILL  FILL_57
timestamp 1490727624
transform 1 0 360 0 -1 290
box -8 -3 16 105
use $$M3_M2  $$M3_M2_153
timestamp 1490727624
transform 1 0 380 0 1 190
box -3 -3 3 3
use NAND2X1  NAND2X1_4
timestamp 1490727624
transform -1 0 392 0 -1 290
box -8 -3 32 105
use LATCH  LATCH_2
timestamp 1490727624
transform 1 0 392 0 -1 290
box -8 -3 64 105
use FILL  FILL_66
timestamp 1490727624
transform 1 0 448 0 -1 290
box -8 -3 16 105
use LATCH  LATCH_3
timestamp 1490727624
transform -1 0 512 0 -1 290
box -8 -3 64 105
use FILL  FILL_67
timestamp 1490727624
transform 1 0 512 0 -1 290
box -8 -3 16 105
use INVX2  INVX2_11
timestamp 1490727624
transform -1 0 536 0 -1 290
box -9 -3 26 105
use FILL  FILL_68
timestamp 1490727624
transform 1 0 536 0 -1 290
box -8 -3 16 105
use FILL  FILL_69
timestamp 1490727624
transform 1 0 544 0 -1 290
box -8 -3 16 105
use AOI21X1  AOI21X1_0
timestamp 1490727624
transform -1 0 584 0 -1 290
box -7 -3 39 105
use FILL  FILL_70
timestamp 1490727624
transform 1 0 584 0 -1 290
box -8 -3 16 105
use FILL  FILL_71
timestamp 1490727624
transform 1 0 592 0 -1 290
box -8 -3 16 105
use FILL  FILL_72
timestamp 1490727624
transform 1 0 600 0 -1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_7
timestamp 1490727624
transform 1 0 608 0 -1 290
box -8 -3 32 105
use FILL  FILL_73
timestamp 1490727624
transform 1 0 632 0 -1 290
box -8 -3 16 105
use NAND3X1  NAND3X1_3
timestamp 1490727624
transform -1 0 672 0 -1 290
box -8 -3 40 105
use FILL  FILL_75
timestamp 1490727624
transform 1 0 672 0 -1 290
box -8 -3 16 105
use NAND3X1  NAND3X1_4
timestamp 1490727624
transform -1 0 712 0 -1 290
box -8 -3 40 105
use FILL  FILL_78
timestamp 1490727624
transform 1 0 712 0 -1 290
box -8 -3 16 105
use FILL  FILL_80
timestamp 1490727624
transform 1 0 720 0 -1 290
box -8 -3 16 105
use INVX2  INVX2_12
timestamp 1490727624
transform -1 0 744 0 -1 290
box -9 -3 26 105
use INVX2  INVX2_13
timestamp 1490727624
transform 1 0 744 0 -1 290
box -9 -3 26 105
use FILL  FILL_86
timestamp 1490727624
transform 1 0 760 0 -1 290
box -8 -3 16 105
use FILL  FILL_87
timestamp 1490727624
transform 1 0 768 0 -1 290
box -8 -3 16 105
use FILL  FILL_88
timestamp 1490727624
transform 1 0 776 0 -1 290
box -8 -3 16 105
use FILL  FILL_89
timestamp 1490727624
transform 1 0 784 0 -1 290
box -8 -3 16 105
use $$M3_M2  $$M3_M2_154
timestamp 1490727624
transform 1 0 804 0 1 190
box -3 -3 3 3
use INVX2  INVX2_14
timestamp 1490727624
transform -1 0 808 0 -1 290
box -9 -3 26 105
use FILL  FILL_90
timestamp 1490727624
transform 1 0 808 0 -1 290
box -8 -3 16 105
use FILL  FILL_91
timestamp 1490727624
transform 1 0 816 0 -1 290
box -8 -3 16 105
use OAI21X1  OAI21X1_5
timestamp 1490727624
transform 1 0 824 0 -1 290
box -8 -3 34 105
use FILL  FILL_92
timestamp 1490727624
transform 1 0 856 0 -1 290
box -8 -3 16 105
use OAI21X1  OAI21X1_6
timestamp 1490727624
transform -1 0 896 0 -1 290
box -8 -3 34 105
use FILL  FILL_99
timestamp 1490727624
transform 1 0 896 0 -1 290
box -8 -3 16 105
use OAI21X1  OAI21X1_7
timestamp 1490727624
transform 1 0 904 0 -1 290
box -8 -3 34 105
use FILL  FILL_100
timestamp 1490727624
transform 1 0 936 0 -1 290
box -8 -3 16 105
use FILL  FILL_105
timestamp 1490727624
transform 1 0 944 0 -1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_8
timestamp 1490727624
transform -1 0 976 0 -1 290
box -8 -3 32 105
use FILL  FILL_106
timestamp 1490727624
transform 1 0 976 0 -1 290
box -8 -3 16 105
use FILL  FILL_107
timestamp 1490727624
transform 1 0 984 0 -1 290
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_7
timestamp 1490727624
transform 1 0 1034 0 1 190
box -7 -2 7 2
use $$M3_M2  $$M3_M2_155
timestamp 1490727624
transform 1 0 4 0 1 160
box -3 -3 3 3
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_8
timestamp 1490727624
transform 1 0 62 0 1 90
box -7 -2 7 2
use FILL  FILL_108
timestamp 1490727624
transform -1 0 88 0 1 90
box -8 -3 16 105
use FILL  FILL_109
timestamp 1490727624
transform -1 0 96 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_156
timestamp 1490727624
transform 1 0 116 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_158
timestamp 1490727624
transform 1 0 116 0 1 140
box -2 -2 2 2
use $$M2_M1  $$M2_M1_160
timestamp 1490727624
transform 1 0 108 0 1 111
box -2 -2 2 2
use $$M3_M2  $$M3_M2_158
timestamp 1490727624
transform 1 0 108 0 1 110
box -3 -3 3 3
use FILL  FILL_110
timestamp 1490727624
transform -1 0 104 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_159
timestamp 1490727624
transform 1 0 124 0 1 133
box -2 -2 2 2
use $$M3_M2  $$M3_M2_157
timestamp 1490727624
transform 1 0 124 0 1 130
box -3 -3 3 3
use NOR2X1  NOR2X1_9
timestamp 1490727624
transform 1 0 104 0 1 90
box -8 -3 32 105
use FILL  FILL_111
timestamp 1490727624
transform -1 0 136 0 1 90
box -8 -3 16 105
use FILL  FILL_112
timestamp 1490727624
transform -1 0 144 0 1 90
box -8 -3 16 105
use FILL  FILL_113
timestamp 1490727624
transform -1 0 152 0 1 90
box -8 -3 16 105
use FILL  FILL_114
timestamp 1490727624
transform -1 0 160 0 1 90
box -8 -3 16 105
use FILL  FILL_115
timestamp 1490727624
transform -1 0 168 0 1 90
box -8 -3 16 105
use FILL  FILL_116
timestamp 1490727624
transform -1 0 176 0 1 90
box -8 -3 16 105
use FILL  FILL_117
timestamp 1490727624
transform -1 0 184 0 1 90
box -8 -3 16 105
use FILL  FILL_118
timestamp 1490727624
transform -1 0 192 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_159
timestamp 1490727624
transform 1 0 204 0 1 170
box -3 -3 3 3
use FILL  FILL_119
timestamp 1490727624
transform -1 0 200 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_161
timestamp 1490727624
transform 1 0 212 0 1 121
box -2 -2 2 2
use $$M3_M2  $$M3_M2_160
timestamp 1490727624
transform 1 0 212 0 1 120
box -3 -3 3 3
use FILL  FILL_120
timestamp 1490727624
transform -1 0 208 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_163
timestamp 1490727624
transform 1 0 244 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_163
timestamp 1490727624
transform 1 0 236 0 1 140
box -3 -3 3 3
use $$M3_M2  $$M3_M2_161
timestamp 1490727624
transform 1 0 220 0 1 110
box -3 -3 3 3
use $$M2_M1  $$M2_M1_162
timestamp 1490727624
transform 1 0 220 0 1 100
box -2 -2 2 2
use INVX2  INVX2_15
timestamp 1490727624
transform 1 0 208 0 1 90
box -9 -3 26 105
use $$M2_M1  $$M2_M1_164
timestamp 1490727624
transform 1 0 236 0 1 133
box -2 -2 2 2
use FILL  FILL_121
timestamp 1490727624
transform -1 0 232 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_162
timestamp 1490727624
transform 1 0 252 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_165
timestamp 1490727624
transform 1 0 244 0 1 120
box -2 -2 2 2
use $$M3_M2  $$M3_M2_164
timestamp 1490727624
transform 1 0 244 0 1 120
box -3 -3 3 3
use $$M2_M1  $$M2_M1_166
timestamp 1490727624
transform 1 0 252 0 1 116
box -2 -2 2 2
use NOR2X1  NOR2X1_10
timestamp 1490727624
transform -1 0 256 0 1 90
box -8 -3 32 105
use $$M3_M2  $$M3_M2_165
timestamp 1490727624
transform 1 0 268 0 1 170
box -3 -3 3 3
use $$M3_M2  $$M3_M2_166
timestamp 1490727624
transform 1 0 284 0 1 170
box -3 -3 3 3
use $$M2_M1  $$M2_M1_167
timestamp 1490727624
transform 1 0 284 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_171
timestamp 1490727624
transform 1 0 268 0 1 127
box -2 -2 2 2
use $$M2_M1  $$M2_M1_169
timestamp 1490727624
transform 1 0 276 0 1 130
box -2 -2 2 2
use $$M3_M2  $$M3_M2_169
timestamp 1490727624
transform 1 0 276 0 1 130
box -3 -3 3 3
use FILL  FILL_122
timestamp 1490727624
transform -1 0 264 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_171
timestamp 1490727624
transform 1 0 292 0 1 110
box -3 -3 3 3
use NAND2X1  NAND2X1_5
timestamp 1490727624
transform 1 0 264 0 1 90
box -8 -3 32 105
use FILL  FILL_123
timestamp 1490727624
transform -1 0 296 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_167
timestamp 1490727624
transform 1 0 324 0 1 160
box -3 -3 3 3
use $$M3_M2  $$M3_M2_168
timestamp 1490727624
transform 1 0 308 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_168
timestamp 1490727624
transform 1 0 316 0 1 137
box -2 -2 2 2
use $$M2_M1  $$M2_M1_170
timestamp 1490727624
transform 1 0 324 0 1 130
box -2 -2 2 2
use $$M2_M1  $$M2_M1_172
timestamp 1490727624
transform 1 0 308 0 1 123
box -2 -2 2 2
use FILL  FILL_124
timestamp 1490727624
transform -1 0 304 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_170
timestamp 1490727624
transform 1 0 324 0 1 120
box -3 -3 3 3
use OAI21X1  OAI21X1_8
timestamp 1490727624
transform 1 0 304 0 1 90
box -8 -3 34 105
use $$M3_M2  $$M3_M2_172
timestamp 1490727624
transform 1 0 348 0 1 170
box -3 -3 3 3
use $$M2_M1  $$M2_M1_173
timestamp 1490727624
transform 1 0 350 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_173
timestamp 1490727624
transform 1 0 350 0 1 150
box -3 -3 3 3
use FILL  FILL_125
timestamp 1490727624
transform -1 0 344 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_174
timestamp 1490727624
transform 1 0 364 0 1 131
box -2 -2 2 2
use $$M2_M1  $$M2_M1_175
timestamp 1490727624
transform 1 0 372 0 1 125
box -2 -2 2 2
use $$M3_M2  $$M3_M2_174
timestamp 1490727624
transform 1 0 372 0 1 110
box -3 -3 3 3
use OAI21X1  OAI21X1_9
timestamp 1490727624
transform -1 0 376 0 1 90
box -8 -3 34 105
use $$M2_M1  $$M2_M1_176
timestamp 1490727624
transform 1 0 388 0 1 139
box -2 -2 2 2
use FILL  FILL_126
timestamp 1490727624
transform -1 0 384 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_175
timestamp 1490727624
transform 1 0 412 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_181
timestamp 1490727624
transform 1 0 420 0 1 143
box -2 -2 2 2
use $$M3_M2  $$M3_M2_179
timestamp 1490727624
transform 1 0 428 0 1 140
box -3 -3 3 3
use $$M3_M2  $$M3_M2_181
timestamp 1490727624
transform 1 0 420 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_182
timestamp 1490727624
transform 1 0 436 0 1 131
box -2 -2 2 2
use $$M3_M2  $$M3_M2_182
timestamp 1490727624
transform 1 0 436 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_178
timestamp 1490727624
transform 1 0 396 0 1 110
box -2 -2 2 2
use $$M3_M2  $$M3_M2_176
timestamp 1490727624
transform 1 0 396 0 1 110
box -3 -3 3 3
use $$M2_M1  $$M2_M1_177
timestamp 1490727624
transform 1 0 412 0 1 111
box -2 -2 2 2
use $$M3_M2  $$M3_M2_177
timestamp 1490727624
transform 1 0 412 0 1 110
box -3 -3 3 3
use $$M2_M1  $$M2_M1_179
timestamp 1490727624
transform 1 0 412 0 1 100
box -2 -2 2 2
use NOR2X1  NOR2X1_11
timestamp 1490727624
transform -1 0 408 0 1 90
box -8 -3 32 105
use FILL  FILL_127
timestamp 1490727624
transform -1 0 416 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_183
timestamp 1490727624
transform 1 0 444 0 1 123
box -2 -2 2 2
use $$M3_M2  $$M3_M2_183
timestamp 1490727624
transform 1 0 444 0 1 100
box -3 -3 3 3
use OAI21X1  OAI21X1_10
timestamp 1490727624
transform -1 0 448 0 1 90
box -8 -3 34 105
use FILL  FILL_128
timestamp 1490727624
transform -1 0 456 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_180
timestamp 1490727624
transform 1 0 468 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_184
timestamp 1490727624
transform 1 0 468 0 1 123
box -2 -2 2 2
use $$M2_M1  $$M2_M1_180
timestamp 1490727624
transform 1 0 484 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_178
timestamp 1490727624
transform 1 0 484 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_185
timestamp 1490727624
transform 1 0 476 0 1 120
box -2 -2 2 2
use $$M3_M2  $$M3_M2_184
timestamp 1490727624
transform 1 0 476 0 1 100
box -3 -3 3 3
use $$M3_M2  $$M3_M2_187
timestamp 1490727624
transform 1 0 468 0 1 90
box -3 -3 3 3
use FILL  FILL_129
timestamp 1490727624
transform -1 0 464 0 1 90
box -8 -3 16 105
use NAND2X1  NAND2X1_6
timestamp 1490727624
transform 1 0 464 0 1 90
box -8 -3 32 105
use $$M2_M1  $$M2_M1_187
timestamp 1490727624
transform 1 0 500 0 1 121
box -2 -2 2 2
use $$M2_M1  $$M2_M1_186
timestamp 1490727624
transform 1 0 508 0 1 160
box -2 -2 2 2
use $$M3_M2  $$M3_M2_185
timestamp 1490727624
transform 1 0 508 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_189
timestamp 1490727624
transform 1 0 516 0 1 110
box -2 -2 2 2
use $$M3_M2  $$M3_M2_186
timestamp 1490727624
transform 1 0 516 0 1 110
box -3 -3 3 3
use $$M3_M2  $$M3_M2_188
timestamp 1490727624
transform 1 0 500 0 1 90
box -3 -3 3 3
use FILL  FILL_130
timestamp 1490727624
transform -1 0 496 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_188
timestamp 1490727624
transform 1 0 524 0 1 121
box -2 -2 2 2
use $$M3_M2  $$M3_M2_189
timestamp 1490727624
transform 1 0 524 0 1 100
box -3 -3 3 3
use INVX2  INVX2_16
timestamp 1490727624
transform 1 0 496 0 1 90
box -9 -3 26 105
use INVX2  INVX2_17
timestamp 1490727624
transform -1 0 528 0 1 90
box -9 -3 26 105
use $$M3_M2  $$M3_M2_190
timestamp 1490727624
transform 1 0 548 0 1 180
box -3 -3 3 3
use $$M3_M2  $$M3_M2_191
timestamp 1490727624
transform 1 0 564 0 1 180
box -3 -3 3 3
use $$M3_M2  $$M3_M2_192
timestamp 1490727624
transform 1 0 556 0 1 170
box -3 -3 3 3
use $$M2_M1  $$M2_M1_190
timestamp 1490727624
transform 1 0 564 0 1 147
box -2 -2 2 2
use $$M2_M1  $$M2_M1_191
timestamp 1490727624
transform 1 0 548 0 1 137
box -2 -2 2 2
use $$M2_M1  $$M2_M1_192
timestamp 1490727624
transform 1 0 540 0 1 123
box -2 -2 2 2
use $$M3_M2  $$M3_M2_193
timestamp 1490727624
transform 1 0 540 0 1 100
box -3 -3 3 3
use FILL  FILL_131
timestamp 1490727624
transform -1 0 536 0 1 90
box -8 -3 16 105
use OAI21X1  OAI21X1_11
timestamp 1490727624
transform 1 0 536 0 1 90
box -8 -3 34 105
use $$M2_M1  $$M2_M1_193
timestamp 1490727624
transform 1 0 588 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_196
timestamp 1490727624
transform 1 0 580 0 1 140
box -2 -2 2 2
use $$M2_M1  $$M2_M1_199
timestamp 1490727624
transform 1 0 596 0 1 137
box -2 -2 2 2
use $$M2_M1  $$M2_M1_197
timestamp 1490727624
transform 1 0 604 0 1 140
box -2 -2 2 2
use $$M2_M1  $$M2_M1_200
timestamp 1490727624
transform 1 0 572 0 1 130
box -2 -2 2 2
use $$M3_M2  $$M3_M2_197
timestamp 1490727624
transform 1 0 596 0 1 120
box -3 -3 3 3
use $$M3_M2  $$M3_M2_198
timestamp 1490727624
transform 1 0 588 0 1 110
box -3 -3 3 3
use $$M3_M2  $$M3_M2_199
timestamp 1490727624
transform 1 0 580 0 1 100
box -3 -3 3 3
use FILL  FILL_132
timestamp 1490727624
transform -1 0 576 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_198
timestamp 1490727624
transform 1 0 612 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_194
timestamp 1490727624
transform 1 0 612 0 1 140
box -3 -3 3 3
use $$M3_M2  $$M3_M2_201
timestamp 1490727624
transform 1 0 604 0 1 90
box -3 -3 3 3
use NAND3X1  NAND3X1_5
timestamp 1490727624
transform -1 0 608 0 1 90
box -8 -3 40 105
use FILL  FILL_133
timestamp 1490727624
transform -1 0 616 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_194
timestamp 1490727624
transform 1 0 644 0 1 180
box -2 -2 2 2
use $$M2_M1  $$M2_M1_195
timestamp 1490727624
transform 1 0 636 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_195
timestamp 1490727624
transform 1 0 628 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_201
timestamp 1490727624
transform 1 0 628 0 1 134
box -2 -2 2 2
use $$M3_M2  $$M3_M2_200
timestamp 1490727624
transform 1 0 636 0 1 120
box -3 -3 3 3
use $$M3_M2  $$M3_M2_196
timestamp 1490727624
transform 1 0 652 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_202
timestamp 1490727624
transform 1 0 652 0 1 130
box -2 -2 2 2
use NAND3X1  NAND3X1_6
timestamp 1490727624
transform 1 0 616 0 1 90
box -8 -3 40 105
use FILL  FILL_134
timestamp 1490727624
transform -1 0 656 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_202
timestamp 1490727624
transform 1 0 676 0 1 180
box -3 -3 3 3
use $$M2_M1  $$M2_M1_203
timestamp 1490727624
transform 1 0 668 0 1 127
box -2 -2 2 2
use $$M3_M2  $$M3_M2_207
timestamp 1490727624
transform 1 0 668 0 1 90
box -3 -3 3 3
use INVX2  INVX2_18
timestamp 1490727624
transform -1 0 672 0 1 90
box -9 -3 26 105
use $$M3_M2  $$M3_M2_205
timestamp 1490727624
transform 1 0 684 0 1 120
box -3 -3 3 3
use $$M2_M1  $$M2_M1_206
timestamp 1490727624
transform 1 0 684 0 1 117
box -2 -2 2 2
use FILL  FILL_135
timestamp 1490727624
transform -1 0 680 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_203
timestamp 1490727624
transform 1 0 700 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_204
timestamp 1490727624
transform 1 0 716 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_204
timestamp 1490727624
transform 1 0 708 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_205
timestamp 1490727624
transform 1 0 700 0 1 133
box -2 -2 2 2
use $$M2_M1  $$M2_M1_207
timestamp 1490727624
transform 1 0 692 0 1 110
box -2 -2 2 2
use $$M3_M2  $$M3_M2_206
timestamp 1490727624
transform 1 0 692 0 1 110
box -3 -3 3 3
use NOR2X1  NOR2X1_12
timestamp 1490727624
transform 1 0 680 0 1 90
box -8 -3 32 105
use FILL  FILL_136
timestamp 1490727624
transform -1 0 712 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_208
timestamp 1490727624
transform 1 0 724 0 1 130
box -2 -2 2 2
use $$M3_M2  $$M3_M2_208
timestamp 1490727624
transform 1 0 724 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_209
timestamp 1490727624
transform 1 0 756 0 1 127
box -2 -2 2 2
use $$M2_M1  $$M2_M1_210
timestamp 1490727624
transform 1 0 740 0 1 110
box -2 -2 2 2
use $$M3_M2  $$M3_M2_209
timestamp 1490727624
transform 1 0 740 0 1 110
box -3 -3 3 3
use NAND2X1  NAND2X1_7
timestamp 1490727624
transform -1 0 736 0 1 90
box -8 -3 32 105
use $$M2_M1  $$M2_M1_211
timestamp 1490727624
transform 1 0 774 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_211
timestamp 1490727624
transform 1 0 774 0 1 180
box -3 -3 3 3
use $$M2_M1  $$M2_M1_212
timestamp 1490727624
transform 1 0 764 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_212
timestamp 1490727624
transform 1 0 788 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_213
timestamp 1490727624
transform 1 0 780 0 1 137
box -2 -2 2 2
use $$M3_M2  $$M3_M2_213
timestamp 1490727624
transform 1 0 780 0 1 130
box -3 -3 3 3
use $$M3_M2  $$M3_M2_214
timestamp 1490727624
transform 1 0 764 0 1 110
box -3 -3 3 3
use $$M3_M2  $$M3_M2_210
timestamp 1490727624
transform 1 0 756 0 1 100
box -3 -3 3 3
use INVX2  INVX2_19
timestamp 1490727624
transform -1 0 752 0 1 90
box -9 -3 26 105
use FILL  FILL_137
timestamp 1490727624
transform -1 0 760 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_214
timestamp 1490727624
transform 1 0 788 0 1 123
box -2 -2 2 2
use OAI21X1  OAI21X1_12
timestamp 1490727624
transform -1 0 792 0 1 90
box -8 -3 34 105
use $$M3_M2  $$M3_M2_215
timestamp 1490727624
transform 1 0 820 0 1 180
box -3 -3 3 3
use $$M2_M1  $$M2_M1_215
timestamp 1490727624
transform 1 0 820 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_216
timestamp 1490727624
transform 1 0 804 0 1 140
box -2 -2 2 2
use FILL  FILL_138
timestamp 1490727624
transform -1 0 800 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_217
timestamp 1490727624
transform 1 0 812 0 1 135
box -2 -2 2 2
use $$M3_M2  $$M3_M2_216
timestamp 1490727624
transform 1 0 812 0 1 110
box -3 -3 3 3
use $$M2_M1  $$M2_M1_218
timestamp 1490727624
transform 1 0 820 0 1 100
box -2 -2 2 2
use $$M3_M2  $$M3_M2_217
timestamp 1490727624
transform 1 0 820 0 1 100
box -3 -3 3 3
use NAND3X1  NAND3X1_7
timestamp 1490727624
transform 1 0 800 0 1 90
box -8 -3 40 105
use $$M3_M2  $$M3_M2_218
timestamp 1490727624
transform 1 0 852 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_219
timestamp 1490727624
transform 1 0 860 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_220
timestamp 1490727624
transform 1 0 844 0 1 140
box -2 -2 2 2
use $$M2_M1  $$M2_M1_221
timestamp 1490727624
transform 1 0 868 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_219
timestamp 1490727624
transform 1 0 868 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_222
timestamp 1490727624
transform 1 0 852 0 1 135
box -2 -2 2 2
use $$M3_M2  $$M3_M2_220
timestamp 1490727624
transform 1 0 844 0 1 130
box -3 -3 3 3
use $$M3_M2  $$M3_M2_221
timestamp 1490727624
transform 1 0 860 0 1 130
box -3 -3 3 3
use FILL  FILL_139
timestamp 1490727624
transform -1 0 840 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_222
timestamp 1490727624
transform 1 0 852 0 1 110
box -3 -3 3 3
use NAND3X1  NAND3X1_8
timestamp 1490727624
transform 1 0 840 0 1 90
box -8 -3 40 105
use $$M2_M1  $$M2_M1_225
timestamp 1490727624
transform 1 0 916 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_225
timestamp 1490727624
transform 1 0 916 0 1 160
box -3 -3 3 3
use $$M3_M2  $$M3_M2_223
timestamp 1490727624
transform 1 0 892 0 1 150
box -3 -3 3 3
use $$M3_M2  $$M3_M2_226
timestamp 1490727624
transform 1 0 908 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_226
timestamp 1490727624
transform 1 0 924 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_223
timestamp 1490727624
transform 1 0 892 0 1 140
box -2 -2 2 2
use $$M2_M1  $$M2_M1_224
timestamp 1490727624
transform 1 0 884 0 1 121
box -2 -2 2 2
use $$M3_M2  $$M3_M2_224
timestamp 1490727624
transform 1 0 884 0 1 120
box -3 -3 3 3
use FILL  FILL_140
timestamp 1490727624
transform -1 0 880 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_227
timestamp 1490727624
transform 1 0 908 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_228
timestamp 1490727624
transform 1 0 900 0 1 90
box -3 -3 3 3
use INVX2  INVX2_20
timestamp 1490727624
transform 1 0 880 0 1 90
box -9 -3 26 105
use FILL  FILL_141
timestamp 1490727624
transform -1 0 904 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_228
timestamp 1490727624
transform 1 0 916 0 1 137
box -2 -2 2 2
use $$M3_M2  $$M3_M2_227
timestamp 1490727624
transform 1 0 924 0 1 130
box -3 -3 3 3
use NAND3X1  NAND3X1_9
timestamp 1490727624
transform 1 0 904 0 1 90
box -8 -3 40 105
use $$M2_M1  $$M2_M1_229
timestamp 1490727624
transform 1 0 961 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_229
timestamp 1490727624
transform 1 0 961 0 1 180
box -3 -3 3 3
use $$M2_M1  $$M2_M1_231
timestamp 1490727624
transform 1 0 948 0 1 117
box -2 -2 2 2
use $$M3_M2  $$M3_M2_233
timestamp 1490727624
transform 1 0 948 0 1 90
box -3 -3 3 3
use FILL  FILL_142
timestamp 1490727624
transform -1 0 944 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_230
timestamp 1490727624
transform 1 0 964 0 1 133
box -2 -2 2 2
use $$M2_M1  $$M2_M1_232
timestamp 1490727624
transform 1 0 980 0 1 130
box -2 -2 2 2
use $$M3_M2  $$M3_M2_231
timestamp 1490727624
transform 1 0 980 0 1 130
box -3 -3 3 3
use $$M3_M2  $$M3_M2_230
timestamp 1490727624
transform 1 0 964 0 1 120
box -3 -3 3 3
use NOR2X1  NOR2X1_13
timestamp 1490727624
transform 1 0 944 0 1 90
box -8 -3 32 105
use FILL  FILL_143
timestamp 1490727624
transform -1 0 976 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_233
timestamp 1490727624
transform 1 0 988 0 1 121
box -2 -2 2 2
use $$M3_M2  $$M3_M2_232
timestamp 1490727624
transform 1 0 988 0 1 120
box -3 -3 3 3
use INVX2  INVX2_21
timestamp 1490727624
transform -1 0 992 0 1 90
box -9 -3 26 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_9
timestamp 1490727624
transform 1 0 1009 0 1 90
box -7 -2 7 2
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_4
timestamp 1490727624
transform 1 0 62 0 1 72
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_5
timestamp 1490727624
transform 1 0 1009 0 1 72
box -7 -7 7 7
use $$M3_M2  $$M3_M2_234
timestamp 1490727624
transform 1 0 4 0 1 60
box -3 -3 3 3
use $$M3_M2  $$M3_M2_235
timestamp 1490727624
transform 1 0 972 0 1 60
box -3 -3 3 3
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_6
timestamp 1490727624
transform 1 0 37 0 1 47
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_7
timestamp 1490727624
transform 1 0 1034 0 1 47
box -7 -7 7 7
<< labels >>
flabel metal3 2 290 2 290 4 FreeSans 26 0 0 0 brnch
flabel metal3 2 170 2 170 4 FreeSans 26 0 0 0 regwrite
flabel metal3 2 60 2 60 4 FreeSans 26 0 0 0 regdst
flabel metal3 2 520 2 520 4 FreeSans 26 0 0 0 iord
flabel metal3 2 400 2 400 4 FreeSans 26 0 0 0 pcwrite
flabel metal2 884 578 884 578 4 FreeSans 26 0 0 0 irwrite[2]
flabel metal2 748 578 748 578 4 FreeSans 26 0 0 0 irwrite[3]
flabel metal2 324 578 324 578 4 FreeSans 26 0 0 0 memwrite
flabel metal2 1028 578 1028 578 4 FreeSans 26 0 0 0 irwrite[1]
flabel metal2 604 578 604 578 4 FreeSans 26 0 0 0 clk
flabel metal2 44 578 44 578 4 FreeSans 26 0 0 0 memtoreg
flabel metal2 188 578 188 578 4 FreeSans 26 0 0 0 alusrca
flabel metal2 468 578 468 578 4 FreeSans 26 0 0 0 reset
flabel metal3 1069 290 1069 290 4 FreeSans 26 0 0 0 aluop[0]
flabel metal3 1069 170 1069 170 4 FreeSans 26 0 0 0 aluop[1]
flabel metal3 1069 400 1069 400 4 FreeSans 26 0 0 0 alusrcb[1]
flabel metal3 1069 520 1069 520 4 FreeSans 26 0 0 0 alusrcb[0]
flabel metal3 1069 60 1069 60 4 FreeSans 26 0 0 0 irwrite[0]
flabel metal2 188 1 188 1 4 FreeSans 26 0 0 0 pcsrc[0]
flabel metal2 884 1 884 1 4 FreeSans 26 0 0 0 op[1]
flabel metal2 1028 1 1028 1 4 FreeSans 26 0 0 0 op[0]
flabel metal2 604 1 604 1 4 FreeSans 26 0 0 0 op[3]
flabel metal2 748 1 748 1 4 FreeSans 26 0 0 0 op[2]
flabel metal2 324 1 324 1 4 FreeSans 26 0 0 0 op[5]
flabel metal2 44 1 44 1 4 FreeSans 26 0 0 0 pcsrc[1]
flabel metal2 468 1 468 1 4 FreeSans 26 0 0 0 op[4]
rlabel metal1 444 71 444 71 1 Gnd!
rlabel metal1 446 45 446 45 1 Vdd!
<< end >>
