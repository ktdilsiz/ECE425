magic
tech scmos
timestamp 1484536911
<< nwell >>
rect 18 40 194 96
<< ntransistor >>
rect 29 7 31 31
rect 37 7 39 13
rect 61 8 63 14
rect 69 8 71 14
rect 85 8 87 14
rect 93 8 95 12
rect 100 8 102 12
rect 109 8 111 14
rect 117 8 119 14
rect 125 8 127 12
rect 132 8 134 12
rect 141 8 143 14
rect 157 8 159 14
rect 165 8 167 14
rect 181 7 183 14
<< ptransistor >>
rect 37 71 39 83
rect 45 77 47 83
rect 61 74 63 83
rect 69 74 71 83
rect 85 77 87 83
rect 93 79 95 83
rect 100 79 102 83
rect 109 74 111 83
rect 117 77 119 83
rect 125 79 127 83
rect 132 79 134 83
rect 141 74 143 83
rect 157 74 159 83
rect 165 74 167 83
rect 181 73 183 83
<< ndiffusion >>
rect 28 7 29 31
rect 31 7 32 31
rect 56 13 61 14
rect 36 7 37 13
rect 39 7 40 13
rect 60 9 61 13
rect 56 8 61 9
rect 63 13 69 14
rect 63 9 64 13
rect 68 9 69 13
rect 63 8 69 9
rect 71 13 76 14
rect 71 9 72 13
rect 71 8 76 9
rect 84 8 85 14
rect 87 8 88 14
rect 104 13 109 14
rect 92 8 93 12
rect 95 8 100 12
rect 102 9 104 12
rect 108 9 109 13
rect 102 8 109 9
rect 111 8 112 14
rect 116 8 117 14
rect 119 8 120 14
rect 136 13 141 14
rect 124 8 125 12
rect 127 8 132 12
rect 134 9 136 12
rect 140 9 141 13
rect 134 8 141 9
rect 143 8 144 14
rect 152 13 157 14
rect 156 9 157 13
rect 152 8 157 9
rect 159 13 165 14
rect 159 9 160 13
rect 164 9 165 13
rect 159 8 165 9
rect 167 8 168 14
rect 176 12 181 14
rect 180 8 181 12
rect 176 7 181 8
rect 183 12 188 14
rect 183 8 184 12
rect 183 7 188 8
<< pdiffusion >>
rect 32 81 37 83
rect 36 72 37 81
rect 32 71 37 72
rect 39 81 45 83
rect 39 72 40 81
rect 44 77 45 81
rect 47 82 52 83
rect 47 78 48 82
rect 47 77 52 78
rect 39 71 44 72
rect 60 74 61 83
rect 63 74 64 83
rect 68 74 69 83
rect 71 74 72 83
rect 80 82 85 83
rect 84 78 85 82
rect 80 77 85 78
rect 87 77 88 83
rect 92 79 93 83
rect 95 79 100 83
rect 102 79 104 83
rect 108 74 109 83
rect 111 74 112 83
rect 116 77 117 83
rect 119 77 120 83
rect 124 79 125 83
rect 127 79 132 83
rect 134 79 136 83
rect 140 74 141 83
rect 143 74 144 83
rect 156 74 157 83
rect 159 74 160 83
rect 164 74 165 83
rect 167 74 168 83
rect 176 82 181 83
rect 180 73 181 82
rect 183 82 188 83
rect 183 73 184 82
<< ndcontact >>
rect 24 7 28 31
rect 32 7 36 31
rect 40 7 44 13
rect 56 9 60 13
rect 64 9 68 13
rect 72 9 76 13
rect 80 8 84 14
rect 88 8 92 14
rect 104 9 108 13
rect 112 8 116 14
rect 120 8 124 14
rect 136 9 140 13
rect 144 8 148 14
rect 152 9 156 13
rect 160 9 164 13
rect 168 8 172 14
rect 176 8 180 12
rect 184 8 188 12
<< pdcontact >>
rect 32 72 36 81
rect 40 72 44 81
rect 48 78 52 82
rect 56 74 60 83
rect 64 74 68 83
rect 72 74 76 83
rect 80 78 84 82
rect 88 77 92 83
rect 104 74 108 83
rect 112 74 116 83
rect 120 77 124 83
rect 136 74 140 83
rect 144 74 148 83
rect 152 74 156 83
rect 160 74 164 83
rect 168 74 172 83
rect 176 73 180 82
rect 184 73 188 82
<< psubstratepcontact >>
rect 24 -2 28 2
rect 32 -2 36 2
rect 40 -2 44 2
rect 48 -2 52 2
rect 56 -2 60 2
rect 64 -2 68 2
rect 72 -2 76 2
rect 80 -2 84 2
rect 88 -2 92 2
rect 96 -2 100 2
rect 104 -2 108 2
rect 112 -2 116 2
rect 120 -2 124 2
rect 128 -2 132 2
rect 136 -2 140 2
rect 144 -2 148 2
rect 152 -2 156 2
rect 160 -2 164 2
rect 168 -2 172 2
rect 176 -2 180 2
rect 184 -2 188 2
<< nsubstratencontact >>
rect 24 88 28 92
rect 32 88 36 92
rect 40 88 44 92
rect 48 88 52 92
rect 56 88 60 92
rect 64 88 68 92
rect 72 88 76 92
rect 80 88 84 92
rect 88 88 92 92
rect 96 88 100 92
rect 104 88 108 92
rect 112 88 116 92
rect 120 88 124 92
rect 128 88 132 92
rect 136 88 140 92
rect 144 88 148 92
rect 152 88 156 92
rect 160 88 164 92
rect 168 88 172 92
rect 176 88 180 92
rect 184 88 188 92
<< polysilicon >>
rect 37 83 39 85
rect 45 83 47 85
rect 61 83 63 85
rect 69 83 71 85
rect 85 83 87 85
rect 93 83 95 85
rect 100 83 102 85
rect 109 83 111 85
rect 117 83 119 85
rect 125 83 127 85
rect 132 83 134 85
rect 141 83 143 85
rect 157 83 159 85
rect 165 83 167 85
rect 181 83 183 85
rect 29 31 31 53
rect 37 47 39 71
rect 45 57 47 77
rect 61 46 63 74
rect 69 57 71 74
rect 85 57 87 77
rect 93 74 95 79
rect 100 67 102 79
rect 100 63 101 67
rect 52 44 63 46
rect 37 13 39 43
rect 61 14 63 44
rect 69 14 71 53
rect 85 45 87 53
rect 85 43 95 45
rect 85 14 87 17
rect 93 12 95 43
rect 100 12 102 63
rect 109 28 111 74
rect 117 57 119 77
rect 125 74 127 79
rect 132 67 134 79
rect 132 63 133 67
rect 120 53 127 55
rect 110 24 111 28
rect 109 14 111 24
rect 117 14 119 17
rect 125 12 127 53
rect 132 12 134 63
rect 141 35 143 74
rect 157 57 159 74
rect 142 31 143 35
rect 141 14 143 31
rect 157 14 159 53
rect 165 33 167 74
rect 165 14 167 29
rect 181 14 183 73
rect 29 5 31 7
rect 37 5 39 7
rect 61 6 63 8
rect 69 6 71 8
rect 85 6 87 8
rect 93 6 95 8
rect 100 6 102 8
rect 109 6 111 8
rect 117 6 119 8
rect 125 6 127 8
rect 132 6 134 8
rect 141 6 143 8
rect 157 6 159 8
rect 165 6 167 8
rect 181 5 183 7
<< polycontact >>
rect 27 53 31 57
rect 44 53 48 57
rect 36 43 40 47
rect 48 43 52 47
rect 92 70 96 74
rect 101 63 105 67
rect 68 53 72 57
rect 84 53 88 57
rect 84 17 88 21
rect 124 70 128 74
rect 133 63 137 67
rect 116 53 120 57
rect 106 24 110 28
rect 116 17 120 21
rect 156 53 160 57
rect 138 31 142 35
rect 177 38 181 42
rect 164 29 168 33
<< metal1 >>
rect 22 92 190 94
rect 22 88 24 92
rect 28 88 32 92
rect 36 88 40 92
rect 44 88 48 92
rect 52 88 56 92
rect 60 88 64 92
rect 68 88 72 92
rect 76 88 80 92
rect 84 88 88 92
rect 92 88 96 92
rect 100 88 104 92
rect 108 88 112 92
rect 116 88 120 92
rect 124 88 128 92
rect 132 88 136 92
rect 140 88 144 92
rect 148 88 152 92
rect 156 88 160 92
rect 164 88 168 92
rect 172 88 176 92
rect 180 88 184 92
rect 188 88 190 92
rect 22 86 190 88
rect 32 81 36 83
rect 32 65 36 72
rect 40 81 44 86
rect 64 83 68 86
rect 104 83 108 86
rect 136 83 140 86
rect 160 83 164 86
rect 40 71 44 72
rect 48 82 52 83
rect 48 71 52 78
rect 80 82 84 83
rect 80 71 84 78
rect 48 67 80 71
rect 112 67 116 74
rect 144 67 148 74
rect 48 65 52 67
rect 32 61 40 65
rect 44 61 52 65
rect 105 63 112 67
rect 137 63 144 67
rect 168 57 172 74
rect 176 82 180 86
rect 184 82 188 83
rect 31 53 44 57
rect 60 53 68 57
rect 72 53 84 57
rect 120 53 156 57
rect 160 53 168 57
rect 56 13 60 53
rect 76 43 96 47
rect 56 8 60 9
rect 64 13 68 14
rect 24 4 28 7
rect 64 4 68 9
rect 72 13 76 43
rect 184 42 188 73
rect 148 38 177 42
rect 124 32 138 35
rect 120 31 138 32
rect 92 24 106 28
rect 132 24 152 28
rect 128 21 132 24
rect 88 17 96 21
rect 120 17 132 21
rect 72 8 76 9
rect 104 13 108 14
rect 104 4 108 9
rect 136 13 140 14
rect 136 4 140 9
rect 152 13 156 24
rect 152 8 156 9
rect 160 13 164 14
rect 160 4 164 9
rect 176 12 180 14
rect 176 4 180 8
rect 184 12 188 38
rect 184 7 188 8
rect 22 2 190 4
rect 22 -2 24 2
rect 28 -2 32 2
rect 36 -2 40 2
rect 44 -2 48 2
rect 52 -2 56 2
rect 60 -2 64 2
rect 68 -2 72 2
rect 76 -2 80 2
rect 84 -2 88 2
rect 92 -2 96 2
rect 100 -2 104 2
rect 108 -2 112 2
rect 116 -2 120 2
rect 124 -2 128 2
rect 132 -2 136 2
rect 140 -2 144 2
rect 148 -2 152 2
rect 156 -2 160 2
rect 164 -2 168 2
rect 172 -2 176 2
rect 180 -2 184 2
rect 188 -2 190 2
rect 22 -4 190 -2
<< m2contact >>
rect 56 74 60 78
rect 72 74 76 78
rect 88 77 92 81
rect 120 77 124 81
rect 152 74 156 78
rect 80 67 84 71
rect 96 70 100 74
rect 128 70 132 74
rect 40 61 44 65
rect 112 63 116 67
rect 144 63 148 67
rect 24 53 27 57
rect 27 53 28 57
rect 56 53 60 57
rect 168 53 172 57
rect 32 43 36 47
rect 48 43 52 47
rect 72 43 76 47
rect 96 43 100 47
rect 40 9 44 13
rect 144 38 148 42
rect 184 38 188 42
rect 120 32 124 36
rect 160 29 164 33
rect 88 24 92 28
rect 128 24 132 28
rect 152 24 156 28
rect 96 17 100 21
rect 80 10 84 14
rect 88 10 92 14
rect 112 10 116 14
rect 120 10 124 14
rect 144 10 148 14
rect 168 10 172 14
<< metal2 >>
rect 40 13 44 61
rect 56 57 60 74
rect 72 47 76 74
rect 80 14 84 67
rect 88 28 92 77
rect 88 14 92 24
rect 96 47 100 70
rect 96 21 100 43
rect 112 14 116 63
rect 120 36 124 77
rect 120 14 124 32
rect 128 28 132 70
rect 144 42 148 63
rect 144 14 148 38
rect 152 28 156 74
rect 168 14 172 53
<< labels >>
rlabel m2contact 26 55 26 55 1 resetb
rlabel metal1 23 90 23 90 3 Vdd!
rlabel metal1 23 0 23 0 3 Gnd!
rlabel m2contact 186 40 186 40 1 q
rlabel m2contact 162 31 162 31 1 ph1
rlabel m2contact 34 45 34 45 1 d
rlabel m2contact 50 45 50 45 1 ph2
rlabel metal1 50 68 50 68 1 masterinb
rlabel metal1 58 32 58 32 1 ph2b
rlabel metal2 170 25 170 25 1 ph1b
rlabel metal1 174 40 174 40 1 slaveb
rlabel metal2 74 63 74 63 1 ph2bb
rlabel metal2 154 33 154 33 1 ph1bb
rlabel metal2 121 37 121 37 1 slave
rlabel metal2 90 36 90 36 1 masterb
rlabel metal2 114 33 114 33 1 master
<< end >>
