magic
tech scmos
timestamp 1492537283
use and2_1x  and2_1x_0
timestamp 1484419738
transform 1 0 5 0 1 4
box -6 -4 34 96
<< end >>
