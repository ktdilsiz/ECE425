magic
tech scmos
timestamp 1487717494
<< nwell >>
rect -6 40 50 96
<< ntransistor >>
rect 5 7 7 28
rect 10 7 12 28
rect 18 7 20 28
rect 23 7 25 28
<< ptransistor >>
rect 5 53 7 83
rect 13 53 15 83
rect 21 53 23 83
rect 29 53 31 83
<< ndiffusion >>
rect 0 27 5 28
rect 4 8 5 27
rect 0 7 5 8
rect 7 7 10 28
rect 12 27 18 28
rect 12 8 13 27
rect 17 8 18 27
rect 12 7 18 8
rect 20 7 23 28
rect 25 27 30 28
rect 25 8 26 27
rect 25 7 30 8
<< pdiffusion >>
rect 0 82 5 83
rect 4 53 5 82
rect 7 82 13 83
rect 7 53 8 82
rect 12 53 13 82
rect 15 82 21 83
rect 15 53 16 82
rect 20 53 21 82
rect 23 82 29 83
rect 23 53 24 82
rect 28 53 29 82
rect 31 76 34 83
rect 31 74 36 76
rect 31 55 32 74
rect 31 53 36 55
<< ndcontact >>
rect 0 8 4 27
rect 13 8 17 27
rect 26 8 30 27
<< pdcontact >>
rect 0 53 4 82
rect 8 53 12 82
rect 16 53 20 82
rect 24 53 28 82
rect 32 55 36 74
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
rect 40 -2 44 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
rect 32 88 36 92
rect 40 88 44 92
<< polysilicon >>
rect 5 83 7 85
rect 13 83 15 85
rect 21 83 23 85
rect 29 83 31 85
rect 5 50 7 53
rect 2 48 7 50
rect 13 49 15 53
rect 2 42 4 48
rect 2 35 4 38
rect 10 47 15 49
rect 10 43 12 47
rect 21 45 23 53
rect 29 52 31 53
rect 29 50 35 52
rect 21 43 26 45
rect 33 43 35 50
rect 24 39 28 43
rect 32 39 36 43
rect 2 33 7 35
rect 5 28 7 33
rect 10 28 12 39
rect 24 36 26 39
rect 18 34 26 36
rect 18 28 20 34
rect 33 31 35 39
rect 23 29 35 31
rect 23 28 25 29
rect 5 5 7 7
rect 10 5 12 7
rect 18 5 20 7
rect 23 5 25 7
<< polycontact >>
rect 0 38 4 42
rect 10 39 14 43
<< metal1 >>
rect -2 92 46 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 32 92
rect 36 88 40 92
rect 44 88 46 92
rect -2 86 46 88
rect 0 82 4 83
rect 8 82 12 86
rect 16 82 20 83
rect 24 82 40 83
rect 28 79 40 82
rect 32 74 36 76
rect 0 50 4 53
rect 16 50 20 53
rect 32 50 36 55
rect 0 46 36 50
rect 14 39 16 43
rect 13 32 40 36
rect 0 27 4 28
rect 0 4 4 8
rect 13 27 17 32
rect 13 7 17 8
rect 26 27 30 28
rect 26 4 30 8
rect -2 2 46 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 40 2
rect 44 -2 46 2
rect -2 -4 46 -2
<< m2contact >>
rect 40 79 44 83
rect 0 38 4 42
rect 16 39 20 43
rect 24 39 28 43
rect 32 39 36 43
rect 40 32 44 36
<< metal2 >>
rect 40 36 44 79
<< labels >>
rlabel m2contact 2 40 2 40 1 b
rlabel m2contact 18 41 18 41 1 a
rlabel m2contact 26 41 26 41 1 c
rlabel m2contact 34 41 34 41 1 d
rlabel m2contact 42 34 42 34 1 y
rlabel metal1 -1 0 -1 0 2 Gnd!
rlabel metal1 -1 90 -1 90 3 Vdd!
<< end >>
