magic
tech scmos
timestamp 1484531287
<< nwell >>
rect -6 40 74 96
<< ntransistor >>
rect 5 7 7 11
rect 13 7 15 11
rect 18 7 20 11
rect 26 7 28 11
rect 43 7 45 11
rect 48 7 50 11
rect 56 7 58 11
rect 61 7 63 11
<< ptransistor >>
rect 5 75 7 83
rect 13 75 15 83
rect 18 75 20 83
rect 26 75 28 83
rect 43 75 45 83
rect 48 75 50 83
rect 56 75 58 83
rect 61 75 63 83
<< ndiffusion >>
rect 4 7 5 11
rect 7 7 8 11
rect 12 7 13 11
rect 15 7 18 11
rect 20 7 21 11
rect 25 7 26 11
rect 28 7 29 11
rect 42 7 43 11
rect 45 7 48 11
rect 50 7 51 11
rect 55 7 56 11
rect 58 7 61 11
rect 63 7 64 11
<< pdiffusion >>
rect 0 81 5 83
rect 4 77 5 81
rect 0 75 5 77
rect 7 81 13 83
rect 7 77 8 81
rect 12 77 13 81
rect 7 75 13 77
rect 15 75 18 83
rect 20 81 26 83
rect 20 77 21 81
rect 25 77 26 81
rect 20 75 26 77
rect 28 81 33 83
rect 28 77 29 81
rect 28 75 33 77
rect 38 81 43 83
rect 42 77 43 81
rect 38 75 43 77
rect 45 75 48 83
rect 50 81 56 83
rect 50 77 51 81
rect 55 77 56 81
rect 50 75 56 77
rect 58 75 61 83
rect 63 81 68 83
rect 63 77 64 81
rect 63 75 68 77
<< ndcontact >>
rect 0 7 4 11
rect 8 7 12 11
rect 21 7 25 11
rect 29 7 33 11
rect 38 7 42 11
rect 51 7 55 11
rect 64 7 68 11
<< pdcontact >>
rect 0 77 4 81
rect 8 77 12 81
rect 21 77 25 81
rect 29 77 33 81
rect 38 77 42 81
rect 51 77 55 81
rect 64 77 68 81
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
rect 40 -2 44 2
rect 48 -2 52 2
rect 56 -2 60 2
rect 64 -2 68 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
rect 32 88 36 92
rect 40 88 44 92
rect 48 88 52 92
rect 56 88 60 92
rect 64 88 68 92
<< polysilicon >>
rect 5 83 7 85
rect 13 83 15 85
rect 18 83 20 85
rect 26 83 28 85
rect 43 83 45 85
rect 48 83 50 85
rect 56 83 58 85
rect 61 83 63 85
rect 5 74 7 75
rect 3 72 7 74
rect 3 51 5 72
rect 13 65 15 75
rect 10 63 15 65
rect 3 14 5 39
rect 10 35 12 63
rect 18 59 20 75
rect 26 71 28 75
rect 10 20 12 31
rect 10 18 15 20
rect 3 12 7 14
rect 5 11 7 12
rect 13 11 15 18
rect 18 11 20 47
rect 26 18 28 67
rect 43 55 45 75
rect 48 74 50 75
rect 56 74 58 75
rect 48 72 58 74
rect 52 47 54 72
rect 61 68 63 75
rect 34 22 36 43
rect 26 11 28 14
rect 43 11 45 25
rect 52 14 54 43
rect 48 12 58 14
rect 48 11 50 12
rect 56 11 58 12
rect 61 11 63 19
rect 5 5 7 7
rect 13 5 15 7
rect 18 5 20 7
rect 26 5 28 7
rect 43 5 45 7
rect 48 5 50 7
rect 56 5 58 7
rect 61 5 63 7
<< polycontact >>
rect 2 47 6 51
rect 2 39 6 43
rect 24 67 28 71
rect 16 55 20 59
rect 17 47 21 51
rect 9 31 13 35
rect 42 51 46 55
rect 60 64 64 68
rect 33 43 37 47
rect 51 43 55 47
rect 42 25 46 29
rect 33 18 37 22
rect 24 14 28 18
rect 60 19 64 23
<< metal1 >>
rect -2 92 70 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 32 92
rect 36 88 40 92
rect 44 88 48 92
rect 52 88 56 92
rect 60 88 64 92
rect 68 88 70 92
rect -2 86 70 88
rect 0 81 4 83
rect 8 81 12 83
rect 8 71 12 77
rect 21 81 25 86
rect 21 75 25 77
rect 29 81 35 83
rect 33 77 35 81
rect 29 75 35 77
rect 8 67 24 71
rect 31 62 35 75
rect 38 81 42 83
rect 38 67 42 77
rect 51 81 55 86
rect 51 75 55 77
rect 64 81 68 83
rect 38 63 40 67
rect 52 64 60 68
rect 38 62 44 63
rect 25 58 35 62
rect 6 47 8 51
rect 12 47 17 51
rect 25 47 29 58
rect 36 51 42 55
rect 25 43 33 47
rect 37 43 51 47
rect 6 39 16 43
rect 25 36 29 43
rect 9 35 29 36
rect 13 32 29 35
rect 28 25 42 29
rect 31 18 33 22
rect 8 14 24 18
rect 8 11 12 14
rect 31 11 35 18
rect 33 7 35 11
rect 38 11 40 15
rect 21 4 25 7
rect 51 4 55 7
rect -2 2 70 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 40 2
rect 44 -2 48 2
rect 52 -2 56 2
rect 60 -2 64 2
rect 68 -2 70 2
rect -2 -4 70 -2
<< m2contact >>
rect 0 77 4 79
rect 0 75 4 77
rect 64 77 68 79
rect 64 75 68 77
rect 40 63 44 67
rect 48 64 52 68
rect 16 55 20 59
rect 8 47 12 51
rect 32 51 36 55
rect 64 53 68 57
rect 16 39 20 43
rect 40 32 44 36
rect 24 25 28 29
rect 0 17 4 21
rect 56 19 60 23
rect 0 7 4 11
rect 40 11 44 15
rect 64 7 68 11
<< metal2 >>
rect 0 21 4 75
rect 16 43 20 55
rect 40 36 44 63
rect 0 11 4 17
rect 40 15 44 32
rect 64 57 68 75
rect 64 11 68 53
<< labels >>
rlabel metal1 -1 0 -1 0 2 Gnd!
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel m2contact 9 49 9 49 1 writeb
rlabel m2contact 18 41 18 41 1 write
rlabel m2contact 50 66 50 66 1 read2b
rlabel m2contact 58 21 58 21 1 read2
rlabel m2contact 26 27 26 27 1 read1
rlabel m2contact 42 34 42 34 1 r1
rlabel m2contact 66 55 66 55 1 r2
rlabel m2contact 2 19 2 19 1 w
rlabel metal1 46 45 46 45 1 data
rlabel metal1 10 69 10 69 1 wt
rlabel m2contact 34 53 34 53 1 read1b
<< end >>
