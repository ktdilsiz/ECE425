magic
tech scmos
timestamp 1484533408
<< metal1 >>
rect 4 318 24 322
rect 33 263 56 267
rect 6 196 46 204
rect 31 152 35 156
rect 31 148 44 152
rect 6 106 46 114
rect 4 98 24 102
rect 22 86 62 94
rect 22 -4 62 4
<< m2contact >>
rect 0 318 4 322
rect 24 318 28 322
rect 56 263 60 267
rect 0 98 4 102
rect 24 98 28 102
<< metal2 >>
rect 24 322 28 386
rect 0 102 4 318
rect 0 2 4 41
rect 0 -2 12 2
rect 16 -2 20 41
rect 24 39 28 98
rect 48 53 52 151
rect 46 52 52 53
rect 46 48 47 52
rect 51 48 52 52
rect 46 47 52 48
rect 32 26 36 41
rect 48 34 52 41
rect 56 39 60 263
rect 64 43 68 151
rect 63 42 69 43
rect 63 38 64 42
rect 68 38 69 42
rect 63 37 69 38
rect 48 30 60 34
rect 32 22 52 26
rect 27 12 33 13
rect 24 8 28 12
rect 32 8 33 12
rect 24 7 33 8
rect 37 12 43 13
rect 37 8 38 12
rect 42 8 43 12
rect 37 7 43 8
rect 24 -2 28 7
rect 38 2 42 7
rect 32 -2 42 2
rect 48 -2 52 22
rect 56 -2 60 30
<< m3contact >>
rect 47 48 51 52
rect 64 38 68 42
rect 28 8 32 12
rect 38 8 42 12
<< metal3 >>
rect 27 52 52 53
rect 27 48 47 52
rect 51 48 52 52
rect 27 47 52 48
rect 27 12 33 47
rect 27 8 28 12
rect 32 8 33 12
rect 27 7 33 8
rect 37 42 69 43
rect 37 38 64 42
rect 68 38 69 42
rect 37 37 69 38
rect 37 12 43 37
rect 37 8 38 12
rect 42 8 43 12
rect 37 7 43 8
use nand5_1x  nand5_1x_0
timestamp 1484533408
transform 1 0 0 0 1 330
box -6 -4 50 96
use nand3_1x  nand3_1x_0
timestamp 1484532417
transform 1 0 8 0 1 220
box -6 -4 34 96
use nand3_1x  nand3_1x_1
timestamp 1484532417
transform 1 0 8 0 1 110
box -6 -4 34 96
use invbuf_4x  invbuf_4x_0
timestamp 1484532969
transform 1 0 40 0 1 110
box -6 -4 34 96
use invbuf_4x  invbuf_4x_1
timestamp 1484532969
transform -1 0 28 0 1 0
box -6 -4 34 96
use invbuf_4x  invbuf_4x_2
timestamp 1484532969
transform -1 0 60 0 1 0
box -6 -4 34 96
<< end >>
