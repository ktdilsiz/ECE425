magic
tech scmos
timestamp 1484534894
<< nwell >>
rect 124 175 125 178
<< metal1 >>
rect 30 856 294 864
rect 348 803 352 807
rect -2 746 294 754
rect -2 662 366 664
rect -2 658 360 662
rect 364 658 366 662
rect -2 656 366 658
rect -2 636 294 644
rect -2 552 366 554
rect -2 548 360 552
rect 364 548 366 552
rect -2 546 366 548
rect -2 526 294 534
rect -2 442 366 444
rect -2 438 360 442
rect 364 438 366 442
rect -2 436 366 438
rect -2 416 294 424
rect -2 332 366 334
rect -2 328 360 332
rect 364 328 366 332
rect -2 326 366 328
rect -2 306 294 314
rect -2 222 366 224
rect -2 218 360 222
rect 364 218 366 222
rect -2 216 366 218
rect -2 196 294 204
rect -2 112 366 114
rect -2 108 360 112
rect 364 108 366 112
rect -2 106 366 108
rect -2 86 294 94
rect 356 33 363 37
rect -2 -4 294 4
<< m2contact >>
rect 344 803 348 807
rect 352 803 356 807
rect 360 768 364 772
rect 360 658 364 662
rect 360 548 364 552
rect 360 438 364 442
rect 360 328 364 332
rect 360 218 364 222
rect 360 108 364 112
rect 352 33 356 37
<< metal2 >>
rect 47 922 53 923
rect 47 918 48 922
rect 52 918 53 922
rect 47 917 53 918
rect 191 922 197 923
rect 191 918 192 922
rect 196 918 197 922
rect 288 918 292 922
rect 320 918 324 922
rect 191 917 197 918
rect 111 852 117 853
rect 111 848 112 852
rect 116 848 117 852
rect 111 847 117 848
rect 143 852 149 853
rect 143 848 144 852
rect 148 848 149 852
rect 143 847 149 848
rect 159 852 165 853
rect 159 848 160 852
rect 164 848 165 852
rect 159 847 165 848
rect 31 842 37 843
rect 31 838 32 842
rect 36 838 37 842
rect 31 837 37 838
rect 95 822 101 823
rect 95 818 96 822
rect 100 818 101 822
rect 95 817 101 818
rect 87 812 93 813
rect 87 808 88 812
rect 92 808 93 812
rect 96 809 100 817
rect 87 807 93 808
rect 112 801 116 847
rect 119 842 125 843
rect 119 838 120 842
rect 124 838 125 842
rect 119 837 125 838
rect 120 832 125 837
rect 144 818 148 847
rect 151 842 157 843
rect 151 838 152 842
rect 156 838 157 842
rect 151 837 157 838
rect 128 803 132 811
rect 127 802 133 803
rect 127 798 128 802
rect 132 798 133 802
rect 127 797 133 798
rect 152 793 156 837
rect 160 803 164 847
rect 167 812 173 813
rect 167 808 168 812
rect 172 808 173 812
rect 167 807 173 808
rect 15 782 21 783
rect 15 778 16 782
rect 20 778 21 782
rect 15 777 21 778
rect 0 673 4 706
rect 16 687 20 777
rect 111 742 117 743
rect 111 738 112 742
rect 116 738 117 742
rect 111 737 117 738
rect 143 742 149 743
rect 143 738 144 742
rect 148 738 149 742
rect 143 737 149 738
rect 159 742 165 743
rect 159 738 160 742
rect 164 738 165 742
rect 159 737 165 738
rect 31 732 37 733
rect 31 728 32 732
rect 36 728 37 732
rect 31 727 37 728
rect 95 712 101 713
rect 95 708 96 712
rect 100 708 101 712
rect 95 707 101 708
rect 87 702 93 703
rect 87 698 88 702
rect 92 698 93 702
rect 96 699 100 707
rect 87 697 93 698
rect 112 691 116 737
rect 119 732 125 733
rect 119 728 120 732
rect 124 728 125 732
rect 119 727 125 728
rect 120 722 125 727
rect 144 708 148 737
rect 151 732 157 733
rect 151 728 152 732
rect 156 728 157 732
rect 151 727 157 728
rect 128 693 132 701
rect 127 692 133 693
rect 127 688 128 692
rect 132 688 133 692
rect 127 687 133 688
rect 152 683 156 727
rect 160 693 164 737
rect 167 702 173 703
rect 167 698 168 702
rect 172 698 173 702
rect 167 697 173 698
rect -1 672 5 673
rect -1 668 0 672
rect 4 668 5 672
rect -1 667 5 668
rect 111 632 117 633
rect 111 628 112 632
rect 116 628 117 632
rect 111 627 117 628
rect 143 632 149 633
rect 143 628 144 632
rect 148 628 149 632
rect 143 627 149 628
rect 159 632 165 633
rect 159 628 160 632
rect 164 628 165 632
rect 159 627 165 628
rect 31 622 37 623
rect 31 618 32 622
rect 36 618 37 622
rect 31 617 37 618
rect 95 602 101 603
rect 95 598 96 602
rect 100 598 101 602
rect 95 597 101 598
rect 87 592 93 593
rect 87 588 88 592
rect 92 588 93 592
rect 96 589 100 597
rect 87 587 93 588
rect 112 581 116 627
rect 119 622 125 623
rect 119 618 120 622
rect 124 618 125 622
rect 119 617 125 618
rect 120 612 125 617
rect 144 598 148 627
rect 151 622 157 623
rect 151 618 152 622
rect 156 618 157 622
rect 151 617 157 618
rect 128 583 132 591
rect 127 582 133 583
rect 127 578 128 582
rect 132 578 133 582
rect 127 577 133 578
rect 152 573 156 617
rect 160 583 164 627
rect 167 592 173 593
rect 167 588 168 592
rect 172 588 173 592
rect 167 587 173 588
rect -1 562 5 563
rect -1 558 0 562
rect 4 558 5 562
rect -1 557 5 558
rect 0 484 4 557
rect 111 522 117 523
rect 111 518 112 522
rect 116 518 117 522
rect 111 517 117 518
rect 143 522 149 523
rect 143 518 144 522
rect 148 518 149 522
rect 143 517 149 518
rect 159 522 165 523
rect 159 518 160 522
rect 164 518 165 522
rect 159 517 165 518
rect 31 512 37 513
rect 31 508 32 512
rect 36 508 37 512
rect 31 507 37 508
rect 95 492 101 493
rect 95 488 96 492
rect 100 488 101 492
rect 95 487 101 488
rect 87 482 93 483
rect 87 478 88 482
rect 92 478 93 482
rect 96 479 100 487
rect 87 477 93 478
rect 112 471 116 517
rect 119 512 125 513
rect 119 508 120 512
rect 124 508 125 512
rect 119 507 125 508
rect 120 502 125 507
rect 144 488 148 517
rect 151 512 157 513
rect 151 508 152 512
rect 156 508 157 512
rect 151 507 157 508
rect 128 473 132 481
rect 127 472 133 473
rect 16 453 20 469
rect 127 468 128 472
rect 132 468 133 472
rect 127 467 133 468
rect 152 463 156 507
rect 160 473 164 517
rect 167 482 173 483
rect 167 478 168 482
rect 172 478 173 482
rect 167 477 173 478
rect 15 452 21 453
rect 15 448 16 452
rect 20 448 21 452
rect 15 447 21 448
rect 111 412 117 413
rect 111 408 112 412
rect 116 408 117 412
rect 111 407 117 408
rect 143 412 149 413
rect 143 408 144 412
rect 148 408 149 412
rect 143 407 149 408
rect 159 412 165 413
rect 159 408 160 412
rect 164 408 165 412
rect 159 407 165 408
rect 31 402 37 403
rect 31 398 32 402
rect 36 398 37 402
rect 31 397 37 398
rect 95 382 101 383
rect 95 378 96 382
rect 100 378 101 382
rect 95 377 101 378
rect 87 372 93 373
rect 87 368 88 372
rect 92 368 93 372
rect 96 369 100 377
rect 87 367 93 368
rect 8 363 12 367
rect 112 361 116 407
rect 119 402 125 403
rect 119 398 120 402
rect 124 398 125 402
rect 119 397 125 398
rect 120 392 125 397
rect 144 378 148 407
rect 151 402 157 403
rect 151 398 152 402
rect 156 398 157 402
rect 151 397 157 398
rect 128 363 132 371
rect 127 362 133 363
rect 127 358 128 362
rect 132 358 133 362
rect 127 357 133 358
rect 152 353 156 397
rect 160 363 164 407
rect 167 372 173 373
rect 167 368 168 372
rect 172 368 173 372
rect 167 367 173 368
rect 15 342 21 343
rect 15 338 16 342
rect 20 338 21 342
rect 15 337 21 338
rect 0 233 4 266
rect 16 247 20 337
rect 111 302 117 303
rect 111 298 112 302
rect 116 298 117 302
rect 111 297 117 298
rect 143 302 149 303
rect 143 298 144 302
rect 148 298 149 302
rect 143 297 149 298
rect 159 302 165 303
rect 159 298 160 302
rect 164 298 165 302
rect 159 297 165 298
rect 31 292 37 293
rect 31 288 32 292
rect 36 288 37 292
rect 95 272 101 273
rect 95 268 96 272
rect 100 268 101 272
rect 95 267 101 268
rect 87 262 93 263
rect 87 258 88 262
rect 92 258 93 262
rect 96 259 100 267
rect 87 257 93 258
rect 112 251 116 297
rect 119 292 125 293
rect 119 288 120 292
rect 124 288 125 292
rect 119 287 125 288
rect 120 285 125 287
rect 120 282 124 285
rect 144 268 148 297
rect 151 292 157 293
rect 151 288 152 292
rect 156 288 157 292
rect 151 287 157 288
rect 128 253 132 261
rect 127 252 133 253
rect 127 248 128 252
rect 132 248 133 252
rect 127 247 133 248
rect 152 243 156 287
rect 160 253 164 297
rect 167 262 173 263
rect 167 258 168 262
rect 172 258 173 262
rect 167 257 173 258
rect -1 232 5 233
rect -1 228 0 232
rect 4 228 5 232
rect -1 227 5 228
rect 111 192 117 193
rect 111 188 112 192
rect 116 188 117 192
rect 111 187 117 188
rect 143 192 149 193
rect 143 188 144 192
rect 148 188 149 192
rect 143 187 149 188
rect 159 192 165 193
rect 159 188 160 192
rect 164 188 165 192
rect 159 187 165 188
rect 95 162 101 163
rect 95 158 96 162
rect 100 158 101 162
rect 95 157 101 158
rect 87 152 93 153
rect 87 148 88 152
rect 92 148 93 152
rect 96 149 100 157
rect 87 147 93 148
rect 112 141 116 187
rect 119 182 125 183
rect 119 178 120 182
rect 124 178 125 182
rect 119 177 125 178
rect 120 175 125 177
rect 120 172 124 175
rect 144 158 148 187
rect 151 182 157 183
rect 151 178 152 182
rect 156 178 157 182
rect 151 177 157 178
rect 128 143 132 151
rect 127 142 133 143
rect 127 138 128 142
rect 132 138 133 142
rect 127 137 133 138
rect 152 133 156 177
rect 160 143 164 187
rect 167 152 173 153
rect 167 148 168 152
rect 172 148 173 152
rect 167 147 173 148
rect 15 122 21 123
rect 15 118 16 122
rect 20 118 21 122
rect 15 117 21 118
rect 0 13 4 46
rect 16 27 20 117
rect 111 82 117 83
rect 111 78 112 82
rect 116 78 117 82
rect 111 77 117 78
rect 143 82 149 83
rect 143 78 144 82
rect 148 78 149 82
rect 143 77 149 78
rect 159 82 165 83
rect 159 78 160 82
rect 164 78 165 82
rect 159 77 165 78
rect 31 72 37 73
rect 31 68 32 72
rect 36 68 37 72
rect 31 67 37 68
rect 95 52 101 53
rect 95 48 96 52
rect 100 48 101 52
rect 95 47 101 48
rect 87 42 93 43
rect 87 38 88 42
rect 92 38 93 42
rect 96 39 100 47
rect 87 37 93 38
rect 112 31 116 77
rect 119 72 125 73
rect 119 68 120 72
rect 124 68 125 72
rect 119 67 125 68
rect 120 65 125 67
rect 120 62 124 65
rect 144 48 148 77
rect 151 72 157 73
rect 151 68 152 72
rect 156 68 157 72
rect 151 67 157 68
rect 128 33 132 41
rect 127 32 133 33
rect 127 28 128 32
rect 132 28 133 32
rect 127 27 133 28
rect 152 23 156 67
rect 160 33 164 77
rect 167 42 173 43
rect 167 38 168 42
rect 172 38 173 42
rect 167 37 173 38
rect 176 23 180 50
rect 192 23 196 917
rect 263 852 269 853
rect 263 848 264 852
rect 268 848 269 852
rect 263 847 269 848
rect 343 852 349 853
rect 343 848 344 852
rect 348 848 349 852
rect 343 847 349 848
rect 264 782 268 847
rect 303 822 309 823
rect 303 818 304 822
rect 308 818 309 822
rect 303 817 309 818
rect 304 805 308 817
rect 344 807 348 847
rect 312 803 316 807
rect 311 802 317 803
rect 311 798 312 802
rect 316 798 317 802
rect 311 797 317 798
rect 263 742 269 743
rect 263 738 264 742
rect 268 738 269 742
rect 263 737 269 738
rect 343 742 349 743
rect 343 738 344 742
rect 348 738 349 742
rect 343 737 349 738
rect 264 672 268 737
rect 303 712 309 713
rect 303 708 304 712
rect 308 708 309 712
rect 344 710 348 737
rect 303 707 309 708
rect 304 695 308 707
rect 312 693 316 697
rect 311 692 317 693
rect 311 688 312 692
rect 316 688 317 692
rect 311 687 317 688
rect 263 632 269 633
rect 263 628 264 632
rect 268 628 269 632
rect 263 627 269 628
rect 343 632 349 633
rect 343 628 344 632
rect 348 628 349 632
rect 343 627 349 628
rect 264 562 268 627
rect 303 602 309 603
rect 303 598 304 602
rect 308 598 309 602
rect 344 600 348 627
rect 303 597 309 598
rect 304 585 308 597
rect 312 583 316 587
rect 311 582 317 583
rect 311 578 312 582
rect 316 578 317 582
rect 311 577 317 578
rect 263 522 269 523
rect 263 518 264 522
rect 268 518 269 522
rect 263 517 269 518
rect 343 522 349 523
rect 343 518 344 522
rect 348 518 349 522
rect 343 517 349 518
rect 264 452 268 517
rect 303 492 309 493
rect 303 488 304 492
rect 308 488 309 492
rect 344 490 348 517
rect 303 487 309 488
rect 304 475 308 487
rect 312 473 316 477
rect 311 472 317 473
rect 311 468 312 472
rect 316 468 317 472
rect 311 467 317 468
rect 263 412 269 413
rect 263 408 264 412
rect 268 408 269 412
rect 263 407 269 408
rect 343 412 349 413
rect 343 408 344 412
rect 348 408 349 412
rect 343 407 349 408
rect 264 342 268 407
rect 303 382 309 383
rect 303 378 304 382
rect 308 378 309 382
rect 344 380 348 407
rect 303 377 309 378
rect 304 365 308 377
rect 312 363 316 367
rect 311 362 317 363
rect 311 358 312 362
rect 316 358 317 362
rect 311 357 317 358
rect 263 302 269 303
rect 263 298 264 302
rect 268 298 269 302
rect 263 297 269 298
rect 343 302 349 303
rect 343 298 344 302
rect 348 298 349 302
rect 343 297 349 298
rect 264 232 268 297
rect 303 272 309 273
rect 303 268 304 272
rect 308 268 309 272
rect 344 270 348 297
rect 303 267 309 268
rect 304 255 308 267
rect 312 253 316 257
rect 311 252 317 253
rect 311 248 312 252
rect 316 248 317 252
rect 311 247 317 248
rect 263 192 269 193
rect 263 188 264 192
rect 268 188 269 192
rect 263 187 269 188
rect 343 192 349 193
rect 343 188 344 192
rect 348 188 349 192
rect 343 187 349 188
rect 264 122 268 187
rect 303 162 309 163
rect 303 158 304 162
rect 308 158 309 162
rect 344 160 348 187
rect 303 157 309 158
rect 304 145 308 157
rect 312 143 316 147
rect 311 142 317 143
rect 311 138 312 142
rect 316 138 317 142
rect 311 137 317 138
rect 263 82 269 83
rect 263 78 264 82
rect 268 78 269 82
rect 263 77 269 78
rect 343 82 349 83
rect 343 78 344 82
rect 348 78 349 82
rect 343 77 349 78
rect 175 22 181 23
rect 175 18 176 22
rect 180 18 181 22
rect 175 17 181 18
rect 191 22 197 23
rect 191 18 192 22
rect 196 18 197 22
rect 191 17 197 18
rect -1 12 5 13
rect 264 12 268 77
rect 303 52 309 53
rect 303 48 304 52
rect 308 48 309 52
rect 344 50 348 77
rect 303 47 309 48
rect 304 35 308 47
rect 352 37 356 803
rect 360 772 364 806
rect 384 783 388 810
rect 383 782 389 783
rect 383 778 384 782
rect 388 778 389 782
rect 383 777 389 778
rect 360 662 364 696
rect 384 673 388 700
rect 383 672 389 673
rect 383 668 384 672
rect 388 668 389 672
rect 383 667 389 668
rect 360 552 364 586
rect 384 563 388 590
rect 383 562 389 563
rect 383 558 384 562
rect 388 558 389 562
rect 383 557 389 558
rect 360 442 364 476
rect 384 453 388 480
rect 383 452 389 453
rect 383 448 384 452
rect 388 448 389 452
rect 383 447 389 448
rect 360 332 364 366
rect 384 343 388 370
rect 383 342 389 343
rect 383 338 384 342
rect 388 338 389 342
rect 383 337 389 338
rect 360 222 364 256
rect 384 233 388 260
rect 383 232 389 233
rect 383 228 384 232
rect 388 228 389 232
rect 383 227 389 228
rect 360 112 364 146
rect 384 123 388 150
rect 383 122 389 123
rect 383 118 384 122
rect 388 118 389 122
rect 383 117 389 118
rect 312 33 316 37
rect 311 32 317 33
rect 311 28 312 32
rect 316 28 317 32
rect 311 27 317 28
rect 384 13 388 40
rect 383 12 389 13
rect -1 8 0 12
rect 4 8 5 12
rect -1 7 5 8
rect 383 8 384 12
rect 388 8 389 12
rect 383 7 389 8
<< m3contact >>
rect 48 918 52 922
rect 192 918 196 922
rect 112 848 116 852
rect 144 848 148 852
rect 160 848 164 852
rect 32 838 36 842
rect 96 818 100 822
rect 88 808 92 812
rect 120 838 124 842
rect 152 838 156 842
rect 128 798 132 802
rect 168 808 172 812
rect 16 778 20 782
rect 112 738 116 742
rect 144 738 148 742
rect 160 738 164 742
rect 32 728 36 732
rect 96 708 100 712
rect 88 698 92 702
rect 120 728 124 732
rect 152 728 156 732
rect 128 688 132 692
rect 168 698 172 702
rect 0 668 4 672
rect 112 628 116 632
rect 144 628 148 632
rect 160 628 164 632
rect 32 618 36 622
rect 96 598 100 602
rect 88 588 92 592
rect 120 618 124 622
rect 152 618 156 622
rect 128 578 132 582
rect 168 588 172 592
rect 0 558 4 562
rect 112 518 116 522
rect 144 518 148 522
rect 160 518 164 522
rect 32 508 36 512
rect 96 488 100 492
rect 88 478 92 482
rect 120 508 124 512
rect 152 508 156 512
rect 128 468 132 472
rect 168 478 172 482
rect 16 448 20 452
rect 112 408 116 412
rect 144 408 148 412
rect 160 408 164 412
rect 32 398 36 402
rect 96 378 100 382
rect 88 368 92 372
rect 120 398 124 402
rect 152 398 156 402
rect 128 358 132 362
rect 168 368 172 372
rect 16 338 20 342
rect 112 298 116 302
rect 144 298 148 302
rect 160 298 164 302
rect 32 288 36 292
rect 96 268 100 272
rect 88 258 92 262
rect 120 288 124 292
rect 152 288 156 292
rect 128 248 132 252
rect 168 258 172 262
rect 0 228 4 232
rect 112 188 116 192
rect 144 188 148 192
rect 160 188 164 192
rect 96 158 100 162
rect 88 148 92 152
rect 120 178 124 182
rect 152 178 156 182
rect 128 138 132 142
rect 168 148 172 152
rect 16 118 20 122
rect 112 78 116 82
rect 144 78 148 82
rect 160 78 164 82
rect 32 68 36 72
rect 96 48 100 52
rect 88 38 92 42
rect 120 68 124 72
rect 152 68 156 72
rect 128 28 132 32
rect 168 38 172 42
rect 264 848 268 852
rect 344 848 348 852
rect 304 818 308 822
rect 312 798 316 802
rect 264 738 268 742
rect 344 738 348 742
rect 304 708 308 712
rect 312 688 316 692
rect 264 628 268 632
rect 344 628 348 632
rect 304 598 308 602
rect 312 578 316 582
rect 264 518 268 522
rect 344 518 348 522
rect 304 488 308 492
rect 312 468 316 472
rect 264 408 268 412
rect 344 408 348 412
rect 304 378 308 382
rect 312 358 316 362
rect 264 298 268 302
rect 344 298 348 302
rect 304 268 308 272
rect 312 248 316 252
rect 264 188 268 192
rect 344 188 348 192
rect 304 158 308 162
rect 312 138 316 142
rect 264 78 268 82
rect 344 78 348 82
rect 176 18 180 22
rect 192 18 196 22
rect 304 48 308 52
rect 384 778 388 782
rect 384 668 388 672
rect 384 558 388 562
rect 384 448 388 452
rect 384 338 388 342
rect 384 228 388 232
rect 384 118 388 122
rect 312 28 316 32
rect 0 8 4 12
rect 384 8 388 12
<< metal3 >>
rect 47 922 197 923
rect 47 918 48 922
rect 52 918 192 922
rect 196 918 197 922
rect 47 917 197 918
rect -17 852 165 853
rect -17 848 112 852
rect 116 848 144 852
rect 148 848 160 852
rect 164 848 165 852
rect -17 847 165 848
rect 263 852 349 853
rect 263 848 264 852
rect 268 848 344 852
rect 348 848 349 852
rect 263 847 349 848
rect -17 842 157 843
rect -17 838 32 842
rect 36 838 120 842
rect 124 838 152 842
rect 156 838 157 842
rect -17 837 157 838
rect 95 822 309 823
rect 95 818 96 822
rect 100 818 304 822
rect 308 818 309 822
rect 95 817 309 818
rect 87 812 173 813
rect 87 808 88 812
rect 92 808 168 812
rect 172 808 173 812
rect 87 807 173 808
rect 127 802 317 803
rect 127 798 128 802
rect 132 798 312 802
rect 316 798 317 802
rect 127 797 317 798
rect -17 782 389 783
rect -17 778 16 782
rect 20 778 384 782
rect 388 778 389 782
rect -17 777 389 778
rect -17 742 165 743
rect -17 738 112 742
rect 116 738 144 742
rect 148 738 160 742
rect 164 738 165 742
rect -17 737 165 738
rect 263 742 349 743
rect 263 738 264 742
rect 268 738 344 742
rect 348 738 349 742
rect 263 737 349 738
rect -17 732 157 733
rect -17 728 32 732
rect 36 728 120 732
rect 124 728 152 732
rect 156 728 157 732
rect -17 727 157 728
rect 95 712 309 713
rect 95 708 96 712
rect 100 708 304 712
rect 308 708 309 712
rect 95 707 309 708
rect 87 702 173 703
rect 87 698 88 702
rect 92 698 168 702
rect 172 698 173 702
rect 87 697 173 698
rect 127 692 317 693
rect 127 688 128 692
rect 132 688 312 692
rect 316 688 317 692
rect 127 687 317 688
rect -17 672 389 673
rect -17 668 0 672
rect 4 668 384 672
rect 388 668 389 672
rect -17 667 389 668
rect -17 632 165 633
rect -17 628 112 632
rect 116 628 144 632
rect 148 628 160 632
rect 164 628 165 632
rect -17 627 165 628
rect 263 632 349 633
rect 263 628 264 632
rect 268 628 344 632
rect 348 628 349 632
rect 263 627 349 628
rect -17 622 157 623
rect -17 618 32 622
rect 36 618 120 622
rect 124 618 152 622
rect 156 618 157 622
rect -17 617 157 618
rect 95 602 309 603
rect 95 598 96 602
rect 100 598 304 602
rect 308 598 309 602
rect 95 597 309 598
rect 87 592 173 593
rect 87 588 88 592
rect 92 588 168 592
rect 172 588 173 592
rect 87 587 173 588
rect 127 582 317 583
rect 127 578 128 582
rect 132 578 312 582
rect 316 578 317 582
rect 127 577 317 578
rect -17 562 389 563
rect -17 558 0 562
rect 4 558 384 562
rect 388 558 389 562
rect -17 557 389 558
rect -17 522 165 523
rect -17 518 112 522
rect 116 518 144 522
rect 148 518 160 522
rect 164 518 165 522
rect -17 517 165 518
rect 263 522 349 523
rect 263 518 264 522
rect 268 518 344 522
rect 348 518 349 522
rect 263 517 349 518
rect -17 512 157 513
rect -17 508 32 512
rect 36 508 120 512
rect 124 508 152 512
rect 156 508 157 512
rect -17 507 157 508
rect 95 492 309 493
rect 95 488 96 492
rect 100 488 304 492
rect 308 488 309 492
rect 95 487 309 488
rect 87 482 173 483
rect 87 478 88 482
rect 92 478 168 482
rect 172 478 173 482
rect 87 477 173 478
rect 127 472 317 473
rect 127 468 128 472
rect 132 468 312 472
rect 316 468 317 472
rect 127 467 317 468
rect -17 452 389 453
rect -17 448 16 452
rect 20 448 384 452
rect 388 448 389 452
rect -17 447 389 448
rect -17 412 165 413
rect -17 408 112 412
rect 116 408 144 412
rect 148 408 160 412
rect 164 408 165 412
rect -17 407 165 408
rect 263 412 349 413
rect 263 408 264 412
rect 268 408 344 412
rect 348 408 349 412
rect 263 407 349 408
rect -17 402 157 403
rect -17 398 32 402
rect 36 398 120 402
rect 124 398 152 402
rect 156 398 157 402
rect -17 397 157 398
rect 95 382 309 383
rect 95 378 96 382
rect 100 378 304 382
rect 308 378 309 382
rect 95 377 309 378
rect 87 372 173 373
rect 87 368 88 372
rect 92 368 168 372
rect 172 368 173 372
rect 87 367 173 368
rect 127 362 317 363
rect 127 358 128 362
rect 132 358 312 362
rect 316 358 317 362
rect 127 357 317 358
rect -17 342 389 343
rect -17 338 16 342
rect 20 338 384 342
rect 388 338 389 342
rect -17 337 389 338
rect -17 302 165 303
rect -17 298 112 302
rect 116 298 144 302
rect 148 298 160 302
rect 164 298 165 302
rect -17 297 165 298
rect 263 302 349 303
rect 263 298 264 302
rect 268 298 344 302
rect 348 298 349 302
rect 263 297 349 298
rect -17 292 157 293
rect -17 288 32 292
rect 36 288 120 292
rect 124 288 152 292
rect 156 288 157 292
rect -17 287 21 288
rect 85 287 157 288
rect 95 272 309 273
rect 95 268 96 272
rect 100 268 304 272
rect 308 268 309 272
rect 95 267 309 268
rect 87 262 173 263
rect 87 258 88 262
rect 92 258 168 262
rect 172 258 173 262
rect 87 257 173 258
rect 127 252 317 253
rect 127 248 128 252
rect 132 248 312 252
rect 316 248 317 252
rect 127 247 317 248
rect -17 232 389 233
rect -17 228 0 232
rect 4 228 384 232
rect 388 228 389 232
rect -17 227 389 228
rect -17 192 165 193
rect -17 188 112 192
rect 116 188 144 192
rect 148 188 160 192
rect 164 188 165 192
rect -17 187 165 188
rect 263 192 349 193
rect 263 188 264 192
rect 268 188 344 192
rect 348 188 349 192
rect 263 187 349 188
rect -17 182 157 183
rect -17 178 120 182
rect 124 178 152 182
rect 156 178 157 182
rect -17 177 157 178
rect 95 162 309 163
rect 95 158 96 162
rect 100 158 304 162
rect 308 158 309 162
rect 95 157 309 158
rect 87 152 173 153
rect 87 148 88 152
rect 92 148 168 152
rect 172 148 173 152
rect 87 147 173 148
rect 127 142 317 143
rect 127 138 128 142
rect 132 138 312 142
rect 316 138 317 142
rect 127 137 317 138
rect -17 122 389 123
rect -17 118 16 122
rect 20 118 384 122
rect 388 118 389 122
rect -17 117 389 118
rect -17 82 165 83
rect -17 78 112 82
rect 116 78 144 82
rect 148 78 160 82
rect 164 78 165 82
rect -17 77 165 78
rect 263 82 349 83
rect 263 78 264 82
rect 268 78 344 82
rect 348 78 349 82
rect 263 77 349 78
rect -17 72 157 73
rect -17 68 32 72
rect 36 68 120 72
rect 124 68 152 72
rect 156 68 157 72
rect -17 67 157 68
rect 95 52 309 53
rect 95 48 96 52
rect 100 48 304 52
rect 308 48 309 52
rect 95 47 309 48
rect 87 42 173 43
rect 87 38 88 42
rect 92 38 168 42
rect 172 38 173 42
rect 87 37 173 38
rect 127 32 317 33
rect 127 28 128 32
rect 132 28 312 32
rect 316 28 317 32
rect 127 27 317 28
rect 175 22 197 23
rect 175 18 176 22
rect 180 18 192 22
rect 196 18 197 22
rect 175 17 197 18
rect -17 12 389 13
rect -17 8 0 12
rect 4 8 384 12
rect 388 8 389 12
rect -17 7 389 8
use yzdetect_8  yzdetect_8_0
timestamp 1484534894
transform 1 0 0 0 1 0
box -8 -4 28 756
use condinv  condinv_0
timestamp 1484534894
transform 1 0 32 0 1 0
box -6 -4 66 976
use and2_1x_8  and2_1x_8_0
timestamp 1484433330
transform 1 0 96 0 1 0
box -6 -4 34 866
use or2_1x_8  or2_1x_8_0
timestamp 1484433330
transform 1 0 128 0 1 0
box -6 -4 34 866
use adder_8  adder_8_0
timestamp 1484427118
transform 1 0 160 0 1 0
box -6 -4 130 866
use mux4_1x_8  mux4_1x_8_0
timestamp 1484532969
transform 1 0 288 0 1 0
box -6 -4 106 976
<< labels >>
rlabel metal3 -15 10 -15 10 3 result_0_
rlabel metal3 -15 69 -15 69 3 b_0_
rlabel metal3 -14 80 -14 80 3 a_0_
rlabel metal3 -14 120 -14 120 3 result_1_
rlabel metal3 -14 180 -14 180 3 b_1_
rlabel metal3 -14 190 -14 190 3 a_1_
rlabel metal3 -14 230 -14 230 3 result_2_
rlabel metal3 -14 290 -14 290 3 b_2_
rlabel metal3 -13 300 -13 300 3 a_2_
rlabel metal3 -13 399 -13 399 3 b_3_
rlabel metal3 -15 510 -15 510 3 b_4_
rlabel metal3 -14 520 -14 520 3 a_4_
rlabel metal3 -14 560 -14 560 3 result_5_
rlabel metal3 -13 620 -13 620 3 b_5_
rlabel metal3 -14 630 -14 630 3 a_5_
rlabel metal3 -14 669 -14 669 3 result_6_
rlabel metal3 -13 730 -13 730 3 b_6_
rlabel metal3 -13 739 -13 739 3 a_6_
rlabel metal3 -14 780 -14 780 3 result_7_
rlabel metal3 -14 839 -14 839 3 b_7_
rlabel metal3 -14 850 -14 850 3 a_7_
rlabel metal3 55 920 55 920 1 alucontrol_2_
rlabel metal1 33 860 33 860 1 Vdd!
rlabel metal1 6 549 6 549 1 Gnd!
rlabel metal1 6 530 6 530 1 Vdd!
rlabel metal1 4 219 4 219 1 Gnd!
rlabel metal1 2 200 2 200 1 Vdd!
rlabel metal1 3 109 3 109 1 Gnd!
rlabel metal1 1 90 1 90 1 Vdd!
rlabel metal1 3 -1 3 -1 1 Gnd!
rlabel metal2 288 918 292 922 1 alucontrol_0_
rlabel metal2 320 918 324 922 1 alucontrol_1_
rlabel metal1 3 310 3 310 1 Vdd!
rlabel metal1 5 330 5 330 1 Gnd!
rlabel metal1 4 419 4 419 1 Vdd!
rlabel metal1 5 440 5 440 1 Gnd!
rlabel metal1 2 640 2 640 1 Vdd!
rlabel metal1 1 659 1 659 1 Gnd!
rlabel metal1 2 749 2 749 1 Vdd!
rlabel metal2 8 363 12 367 1 zero
rlabel metal3 -13 340 -13 340 3 result_3_
rlabel metal3 -14 450 -14 450 3 result_4_
rlabel metal3 -14 410 -14 410 3 a_3_
<< end >>
