magic
tech scmos
timestamp 1485892876
<< nwell >>
rect -63 8 41 36
rect -19 -10 9 8
<< ntransistor >>
rect -47 -7 -39 -5
rect 16 -11 20 -9
rect -47 -15 -39 -13
<< ptransistor >>
rect -47 21 -31 23
rect 15 21 31 23
rect -13 7 3 9
<< ndiffusion >>
rect -47 -5 -39 -4
rect -47 -13 -39 -7
rect 16 -9 20 -4
rect -47 -16 -39 -15
rect 16 -16 20 -11
<< pdiffusion >>
rect -47 23 -31 24
rect 15 23 31 24
rect -47 20 -31 21
rect 15 20 31 21
rect -13 9 3 14
rect -13 2 3 7
<< ndcontact >>
rect -47 -4 -39 2
rect 16 -4 20 2
rect -47 -22 -39 -16
rect 16 -22 20 -16
<< pdcontact >>
rect -47 24 -31 30
rect 15 24 31 30
rect -47 14 -31 20
rect -13 14 3 20
rect 15 14 31 20
rect -13 -4 3 2
<< polysilicon >>
rect -54 21 -47 23
rect -31 21 -28 23
rect -25 21 15 23
rect 31 21 34 23
rect -54 1 -52 21
rect -58 -1 -52 1
rect -54 -5 -52 -1
rect -54 -7 -47 -5
rect -39 -7 -37 -5
rect -25 -13 -23 21
rect -15 7 -13 9
rect 3 7 10 9
rect 8 -9 10 7
rect 8 -11 16 -9
rect 20 -11 27 -9
rect -57 -15 -47 -13
rect -39 -15 -23 -13
<< polycontact >>
rect -62 -2 -58 2
rect -61 -16 -57 -12
rect -19 6 -15 10
<< metal1 >>
rect -51 24 -47 30
rect -31 24 15 30
rect 31 24 34 30
rect -51 14 -47 20
rect -31 14 -13 20
rect 3 14 15 20
rect 31 14 34 20
rect -59 6 -19 10
rect -65 -2 -62 2
rect -51 -4 -47 2
rect -39 -4 -13 2
rect 3 -4 16 2
rect 20 -4 30 2
rect -65 -16 -61 -12
rect -51 -22 -47 -16
rect -39 -22 16 -16
rect 20 -22 30 -16
<< labels >>
rlabel metal1 -49 27 -49 27 5 Vdd!
rlabel metal1 -64 -14 -64 -14 1 B
rlabel metal1 -57 8 -57 8 1 C
rlabel metal1 -64 0 -64 0 3 A
rlabel metal1 26 -19 26 -19 8 Gnd!
rlabel metal1 27 -1 27 -1 7 Y
<< end >>
