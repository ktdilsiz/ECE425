magic
tech scmos
timestamp 1494344105
<< metal1 >>
rect 1003 3996 1351 3997
rect 1003 3992 1346 3996
rect 1350 3992 1351 3996
rect 1003 3991 1351 3992
rect 1003 1257 1009 3991
rect 1012 3984 1646 3988
rect 1012 1354 1016 3984
rect 1019 3977 1946 3981
rect 1019 1464 1023 3977
rect 1026 3970 2246 3974
rect 1026 1571 1030 3970
rect 1033 3963 2546 3967
rect 2550 3963 2551 3967
rect 1033 1684 1037 3963
rect 1040 3957 2846 3960
rect 1040 3956 2850 3957
rect 1040 1791 1044 3956
rect 1134 3879 1233 3886
rect 1383 3881 1474 3886
rect 1134 3875 1239 3879
rect 1134 3866 1253 3875
rect 1383 3870 1491 3881
rect 1134 3857 1263 3866
rect 1383 3857 1507 3870
rect 1134 3852 1277 3857
rect 1134 3625 1168 3852
rect 1199 3851 1277 3852
rect 1383 3852 1524 3857
rect 1199 3845 1286 3851
rect 1205 3841 1286 3845
rect 1219 3840 1286 3841
rect 1219 3834 1297 3840
rect 1219 3832 1309 3834
rect 1229 3823 1309 3832
rect 1243 3817 1309 3823
rect 1252 3806 1317 3817
rect 1263 3800 1317 3806
rect 1272 3783 1317 3800
rect 1283 3745 1317 3783
rect 1383 3751 1417 3852
rect 1440 3847 1524 3852
rect 1457 3840 1524 3847
rect 1617 3855 1816 3889
rect 1935 3888 1991 3895
rect 1935 3880 1998 3888
rect 1919 3874 1998 3880
rect 2097 3885 2152 3893
rect 2097 3877 2161 3885
rect 2338 3878 2382 3889
rect 2642 3879 2779 3892
rect 2839 3882 2894 3890
rect 2642 3878 2791 3879
rect 1919 3867 2013 3874
rect 1457 3836 1537 3840
rect 1473 3823 1537 3836
rect 1490 3806 1537 3823
rect 1503 3781 1537 3806
rect 1498 3774 1537 3781
rect 1481 3764 1537 3774
rect 1442 3751 1537 3764
rect 1383 3747 1537 3751
rect 1617 3761 1651 3855
rect 1782 3846 1816 3855
rect 1903 3865 2013 3867
rect 1903 3853 2017 3865
rect 2097 3863 2174 3877
rect 2327 3863 2382 3878
rect 1903 3846 2024 3853
rect 1903 3834 1953 3846
rect 1964 3841 2024 3846
rect 2097 3848 2185 3863
rect 2309 3848 2382 3863
rect 2097 3843 2195 3848
rect 1964 3840 2035 3841
rect 1882 3833 1953 3834
rect 1882 3807 1937 3833
rect 1979 3831 2035 3840
rect 1983 3823 2035 3831
rect 1983 3819 2045 3823
rect 1990 3807 2045 3819
rect 1868 3800 1937 3807
rect 2001 3803 2045 3807
rect 1868 3789 1916 3800
rect 2001 3790 2053 3803
rect 2001 3789 2061 3790
rect 1858 3776 1916 3789
rect 1841 3773 1916 3776
rect 2011 3778 2061 3789
rect 1383 3745 1532 3747
rect 1283 3711 1318 3745
rect 1382 3740 1532 3745
rect 1382 3730 1515 3740
rect 1382 3717 1476 3730
rect 1617 3727 1709 3761
rect 1841 3755 1902 3773
rect 2011 3769 2072 3778
rect 2019 3756 2072 3769
rect 1841 3742 1892 3755
rect 2027 3744 2072 3756
rect 1382 3712 1464 3717
rect 1382 3711 1473 3712
rect 1283 3690 1317 3711
rect 1276 3681 1317 3690
rect 1265 3669 1317 3681
rect 1251 3656 1317 3669
rect 1251 3654 1310 3656
rect 1235 3647 1310 3654
rect 1235 3644 1299 3647
rect 1229 3635 1299 3644
rect 1210 3625 1285 3635
rect 1134 3620 1285 3625
rect 1134 3610 1269 3620
rect 1134 3601 1263 3610
rect 1134 3591 1244 3601
rect 1383 3585 1417 3711
rect 1420 3703 1473 3711
rect 1420 3695 1483 3703
rect 1430 3688 1483 3695
rect 1430 3678 1493 3688
rect 1439 3675 1493 3678
rect 1439 3669 1510 3675
rect 1449 3666 1510 3669
rect 1449 3655 1527 3666
rect 1449 3654 1539 3655
rect 1459 3645 1539 3654
rect 1459 3641 1552 3645
rect 1476 3634 1552 3641
rect 1476 3632 1565 3634
rect 1493 3624 1565 3632
rect 1617 3624 1651 3727
rect 1841 3724 1875 3742
rect 2038 3724 2072 3744
rect 1841 3690 2072 3724
rect 1779 3624 1813 3629
rect 1493 3621 1568 3624
rect 1505 3611 1568 3621
rect 1518 3600 1568 3611
rect 1531 3590 1568 3600
rect 1615 3590 1813 3624
rect 1841 3624 1875 3690
rect 1841 3590 1876 3624
rect 2038 3620 2072 3690
rect 2038 3586 2073 3620
rect 2097 3586 2131 3843
rect 2140 3836 2195 3843
rect 2140 3829 2203 3836
rect 2297 3832 2382 3848
rect 2594 3861 2791 3878
rect 2839 3874 2903 3882
rect 3080 3875 3124 3886
rect 3240 3883 3296 3890
rect 3240 3875 3303 3883
rect 2594 3858 2797 3861
rect 2594 3845 2676 3858
rect 2716 3849 2797 3858
rect 2745 3845 2797 3849
rect 2151 3821 2203 3829
rect 2280 3829 2382 3832
rect 2151 3814 2211 3821
rect 2280 3816 2343 3829
rect 2161 3809 2211 3814
rect 2269 3814 2343 3816
rect 2161 3802 2218 3809
rect 2169 3799 2218 3802
rect 2269 3799 2331 3814
rect 2169 3787 2232 3799
rect 2177 3781 2232 3787
rect 2249 3798 2331 3799
rect 2249 3782 2314 3798
rect 2177 3777 2241 3781
rect 2249 3777 2303 3782
rect 2177 3775 2303 3777
rect 2184 3765 2303 3775
rect 2198 3747 2283 3765
rect 2207 3743 2283 3747
rect 2207 3742 2275 3743
rect 2215 3727 2275 3742
rect 2348 3620 2382 3829
rect 2583 3844 2676 3845
rect 2583 3811 2628 3844
rect 2757 3827 2797 3845
rect 2763 3811 2797 3827
rect 2839 3860 2916 3874
rect 3069 3860 3124 3875
rect 3224 3869 3303 3875
rect 3224 3862 3318 3869
rect 2839 3845 2927 3860
rect 3051 3845 3124 3860
rect 2839 3840 2937 3845
rect 2583 3782 2617 3811
rect 2583 3772 2630 3782
rect 2583 3755 2664 3772
rect 2583 3748 2703 3755
rect 2596 3738 2703 3748
rect 2630 3733 2703 3738
rect 2630 3721 2756 3733
rect 2669 3699 2788 3721
rect 2722 3687 2788 3699
rect 2740 3659 2788 3687
rect 2574 3652 2608 3658
rect 2740 3655 2774 3659
rect 2574 3635 2613 3652
rect 2728 3644 2774 3655
rect 2574 3623 2627 3635
rect 2719 3629 2774 3644
rect 2574 3620 2635 3623
rect 2702 3621 2774 3629
rect 2702 3620 2762 3621
rect 2348 3609 2383 3620
rect 2574 3618 2762 3620
rect 2346 3586 2383 3609
rect 2579 3610 2762 3618
rect 2579 3601 2753 3610
rect 2593 3595 2753 3601
rect 2593 3589 2736 3595
rect 2601 3586 2736 3589
rect 2038 3585 2072 3586
rect 2839 3583 2873 3840
rect 2882 3833 2937 3840
rect 2882 3826 2945 3833
rect 3039 3829 3124 3845
rect 3208 3860 3318 3862
rect 3208 3848 3322 3860
rect 3208 3841 3329 3848
rect 3208 3829 3258 3841
rect 3269 3836 3329 3841
rect 3269 3835 3340 3836
rect 2893 3818 2945 3826
rect 3022 3826 3124 3829
rect 2893 3811 2953 3818
rect 3022 3813 3085 3826
rect 2903 3806 2953 3811
rect 3011 3811 3085 3813
rect 2903 3799 2960 3806
rect 2911 3796 2960 3799
rect 3011 3796 3073 3811
rect 2911 3784 2974 3796
rect 2919 3778 2974 3784
rect 2991 3795 3073 3796
rect 2991 3779 3056 3795
rect 2919 3774 2983 3778
rect 2991 3774 3045 3779
rect 2919 3772 3045 3774
rect 2926 3762 3045 3772
rect 2940 3744 3025 3762
rect 2949 3740 3025 3744
rect 2949 3739 3017 3740
rect 2957 3724 3017 3739
rect 3090 3617 3124 3826
rect 3187 3828 3258 3829
rect 3187 3802 3242 3828
rect 3284 3826 3340 3835
rect 3288 3818 3340 3826
rect 3288 3814 3350 3818
rect 3295 3802 3350 3814
rect 3173 3795 3242 3802
rect 3306 3798 3350 3802
rect 3173 3784 3221 3795
rect 3306 3785 3358 3798
rect 3306 3784 3366 3785
rect 3163 3771 3221 3784
rect 3146 3768 3221 3771
rect 3316 3773 3366 3784
rect 3146 3750 3207 3768
rect 3316 3764 3377 3773
rect 3324 3751 3377 3764
rect 3146 3737 3197 3750
rect 3332 3739 3377 3751
rect 3146 3719 3180 3737
rect 3343 3719 3377 3739
rect 3146 3685 3377 3719
rect 3146 3619 3180 3685
rect 3090 3606 3125 3617
rect 3088 3583 3125 3606
rect 3146 3585 3181 3619
rect 3343 3585 3377 3685
rect 3419 3619 3453 3893
rect 3671 3619 3705 3904
rect 3961 3850 4007 3851
rect 3965 3846 4007 3850
rect 3961 3845 4007 3846
rect 3418 3585 3643 3619
rect 3671 3585 3879 3619
rect 3968 3550 4006 3551
rect 3972 3546 4006 3550
rect 3968 3544 4006 3546
rect 2784 3386 2872 3406
rect 2905 3404 2925 3518
rect 2972 3439 2983 3442
rect 2963 3435 2983 3439
rect 2956 3430 2983 3435
rect 2949 3428 2983 3430
rect 3024 3433 3038 3446
rect 2949 3424 2978 3428
rect 2949 3422 2967 3424
rect 2943 3419 2967 3422
rect 2943 3417 2960 3419
rect 2938 3411 2960 3417
rect 3024 3416 3037 3433
rect 2938 3409 2954 3411
rect 2929 3406 2954 3409
rect 2929 3404 2949 3406
rect 2905 3400 2949 3404
rect 3007 3403 3050 3416
rect 2905 3397 2940 3400
rect 2905 3387 2947 3397
rect 2905 3384 2958 3387
rect 2905 3329 2925 3384
rect 2934 3375 2964 3384
rect 2934 3374 2973 3375
rect 2945 3371 2973 3374
rect 2951 3366 2973 3371
rect 2951 3362 2981 3366
rect 2960 3356 2981 3362
rect 2960 3353 2988 3356
rect 2968 3345 2988 3353
rect 3024 3351 3037 3403
rect 3142 3402 3155 3519
rect 3182 3431 3195 3433
rect 3178 3418 3201 3431
rect 3182 3417 3195 3418
rect 3102 3396 3155 3402
rect 3093 3389 3155 3396
rect 3093 3383 3115 3389
rect 3093 3359 3106 3383
rect 3093 3351 3121 3359
rect 2968 3343 2994 3345
rect 2975 3332 2994 3343
rect 2981 3326 2994 3332
rect 3024 3344 3046 3351
rect 3060 3346 3076 3349
rect 3093 3346 3128 3351
rect 3142 3346 3155 3389
rect 3058 3344 3076 3346
rect 3024 3336 3076 3344
rect 3108 3338 3155 3346
rect 3024 3333 3073 3336
rect 3115 3333 3155 3338
rect 3182 3333 3195 3407
rect 3223 3352 3236 3519
rect 3402 3430 3415 3431
rect 3402 3429 3419 3430
rect 3314 3422 3352 3424
rect 3314 3419 3358 3422
rect 3300 3411 3358 3419
rect 3395 3417 3419 3429
rect 3395 3416 3417 3417
rect 3402 3415 3417 3416
rect 3450 3411 3525 3424
rect 3300 3406 3327 3411
rect 3345 3406 3358 3411
rect 3512 3407 3525 3411
rect 3300 3394 3313 3406
rect 3300 3383 3322 3394
rect 3300 3381 3352 3383
rect 3309 3379 3352 3381
rect 3309 3370 3361 3379
rect 3339 3366 3361 3370
rect 3348 3360 3361 3366
rect 3223 3347 3247 3352
rect 3261 3347 3274 3351
rect 3223 3334 3274 3347
rect 3298 3350 3311 3352
rect 3339 3351 3361 3360
rect 3298 3348 3318 3350
rect 3298 3347 3322 3348
rect 3334 3347 3361 3351
rect 3298 3338 3352 3347
rect 3298 3337 3347 3338
rect 3305 3335 3347 3337
rect 3402 3335 3415 3403
rect 3507 3395 3525 3407
rect 3500 3394 3525 3395
rect 3500 3388 3520 3394
rect 3493 3382 3520 3388
rect 3493 3379 3513 3382
rect 3478 3375 3513 3379
rect 3478 3373 3506 3375
rect 3469 3366 3506 3373
rect 3469 3365 3491 3366
rect 3461 3360 3491 3365
rect 3461 3356 3482 3360
rect 3454 3352 3482 3356
rect 3454 3351 3474 3352
rect 3450 3348 3474 3351
rect 3450 3335 3523 3348
rect 3309 3334 3347 3335
rect 3223 3333 3236 3334
rect 3024 3331 3071 3333
rect 2904 3275 2960 3276
rect 2904 3271 3965 3275
rect 2904 3267 3961 3271
rect 2904 3262 3965 3267
rect 2904 3261 2960 3262
rect 2904 3212 2916 3261
rect 1105 3200 1208 3207
rect 1105 3176 1109 3200
rect 1067 3086 1074 3094
rect 1067 2991 1071 3086
rect 1119 3080 1124 3200
rect 2205 3198 2916 3212
rect 2920 3237 2935 3239
rect 2920 3235 2941 3237
rect 2920 3230 2935 3235
rect 2940 3230 2941 3235
rect 2920 3228 2941 3230
rect 2920 3185 2935 3228
rect 2176 3173 2935 3185
rect 1104 3074 1124 3080
rect 2920 3030 2935 3173
rect 2929 3021 2935 3030
rect 2945 2998 2960 3261
rect 2964 3235 3972 3237
rect 2964 3230 2965 3235
rect 2970 3231 3968 3235
rect 2970 3230 3972 3231
rect 2964 3228 3972 3230
rect 3815 3134 3965 3135
rect 3815 3130 3961 3134
rect 3815 3127 3965 3130
rect 3815 3043 3972 3045
rect 3815 3039 3968 3043
rect 3815 3037 3972 3039
rect 3815 3003 3965 3005
rect 3815 2999 3961 3003
rect 3815 2997 3965 2999
rect 1067 2990 1074 2991
rect 1067 2989 1076 2990
rect 1067 2985 1069 2989
rect 1073 2985 1076 2989
rect 1067 2984 1076 2985
rect 1067 2983 1074 2984
rect 3815 2913 3972 2915
rect 3815 2909 3968 2913
rect 3815 2907 3972 2909
rect 3815 2873 3965 2875
rect 3815 2869 3961 2873
rect 3815 2867 3965 2869
rect 3815 2783 3972 2785
rect 3815 2779 3968 2783
rect 3815 2777 3972 2779
rect 3815 2743 3965 2745
rect 3815 2739 3961 2743
rect 3815 2737 3965 2739
rect 3815 2654 3972 2655
rect 3815 2650 3968 2654
rect 3815 2647 3972 2650
rect 3910 2484 3965 2486
rect 3910 2480 3961 2484
rect 3910 2478 3965 2480
rect 3958 2394 3972 2396
rect 3958 2390 3968 2394
rect 3958 2388 3972 2390
rect 3910 2375 3965 2376
rect 3910 2371 3961 2375
rect 3910 2368 3965 2371
rect 3958 2284 3972 2286
rect 3958 2280 3968 2284
rect 3958 2278 3972 2280
rect 3910 2264 3965 2266
rect 3910 2260 3961 2264
rect 3910 2258 3965 2260
rect 3958 2174 3972 2176
rect 3958 2170 3968 2174
rect 3958 2168 3972 2170
rect 3910 2155 3965 2156
rect 3910 2151 3961 2155
rect 3910 2148 3965 2151
rect 3958 2064 3972 2066
rect 3958 2060 3968 2064
rect 3958 2058 3972 2060
rect 3910 2044 3965 2046
rect 3910 2040 3961 2044
rect 3910 2038 3965 2040
rect 3958 1954 3972 1956
rect 3958 1950 3968 1954
rect 3958 1948 3972 1950
rect 3910 1934 3965 1936
rect 3910 1930 3961 1934
rect 3910 1928 3965 1930
rect 1180 1900 1182 1904
rect 1186 1900 1209 1904
rect 3958 1844 3972 1846
rect 3958 1840 3968 1844
rect 3958 1838 3972 1840
rect 3910 1824 3965 1826
rect 3910 1820 3961 1824
rect 3910 1818 3965 1820
rect 1040 1790 1211 1791
rect 1040 1787 1215 1790
rect 3958 1734 3972 1736
rect 3958 1730 3968 1734
rect 3958 1728 3972 1730
rect 3910 1715 3965 1716
rect 3910 1711 3961 1715
rect 3910 1708 3965 1711
rect 1033 1680 1211 1684
rect 3958 1624 3972 1626
rect 3958 1620 3968 1624
rect 3958 1618 3972 1620
rect 3910 1604 3965 1606
rect 3910 1600 3961 1604
rect 3910 1598 3965 1600
rect 1203 1571 1213 1573
rect 1026 1570 1213 1571
rect 1026 1569 1217 1570
rect 1026 1567 1207 1569
rect 3958 1514 3972 1516
rect 3958 1510 3968 1514
rect 3958 1508 3972 1510
rect 3910 1494 3965 1496
rect 3910 1490 3961 1494
rect 3910 1488 3965 1490
rect 1019 1460 1203 1464
rect 3958 1404 3972 1406
rect 3958 1400 3968 1404
rect 3958 1398 3972 1400
rect 3910 1384 3965 1386
rect 3910 1380 3961 1384
rect 3910 1378 3965 1380
rect 1012 1350 1204 1354
rect 1208 1350 1212 1354
rect 3958 1294 3972 1296
rect 3958 1290 3968 1294
rect 3958 1288 3972 1290
rect 3910 1274 3965 1276
rect 3910 1270 3961 1274
rect 3910 1268 3965 1270
rect 1003 1251 1042 1257
rect 1036 1245 1042 1251
rect 3958 1184 3972 1186
rect 3958 1180 3968 1184
rect 3958 1178 3972 1180
<< m2contact >>
rect 1346 3992 1350 3996
rect 1646 3984 1650 3988
rect 1946 3977 1950 3981
rect 2246 3970 2250 3974
rect 2546 3963 2550 3967
rect 2846 3957 2850 3961
rect 3961 3846 3965 3850
rect 3968 3546 3972 3550
rect 3961 3267 3965 3271
rect 2935 3230 2940 3235
rect 2920 3021 2929 3030
rect 2965 3230 2970 3235
rect 3968 3231 3972 3235
rect 3961 3130 3965 3134
rect 3968 3039 3972 3043
rect 3961 2999 3965 3003
rect 1069 2985 1073 2989
rect 3968 2909 3972 2913
rect 3961 2869 3965 2873
rect 3968 2779 3972 2783
rect 3961 2739 3965 2743
rect 3968 2650 3972 2654
rect 3961 2480 3965 2484
rect 3968 2390 3972 2394
rect 3961 2371 3965 2375
rect 3968 2280 3972 2284
rect 3961 2260 3965 2264
rect 3968 2170 3972 2174
rect 3961 2151 3965 2155
rect 3968 2060 3972 2064
rect 3961 2040 3965 2044
rect 3968 1950 3972 1954
rect 3961 1930 3965 1934
rect 1182 1900 1186 1904
rect 1209 1900 1213 1904
rect 3968 1840 3972 1844
rect 3961 1820 3965 1824
rect 1211 1790 1215 1794
rect 3968 1730 3972 1734
rect 3961 1711 3965 1715
rect 1211 1680 1215 1684
rect 3968 1620 3972 1624
rect 3961 1600 3965 1604
rect 1213 1570 1217 1574
rect 3968 1510 3972 1514
rect 3961 1490 3965 1494
rect 1203 1460 1207 1464
rect 3968 1400 3972 1404
rect 3961 1380 3965 1384
rect 1204 1350 1208 1354
rect 3968 1290 3972 1294
rect 3961 1270 3965 1274
rect 1036 1239 1042 1245
rect 3968 1180 3972 1184
<< metal2 >>
rect 1259 3998 1263 4000
rect 1345 3996 1351 4010
rect 1345 3992 1346 3996
rect 1350 3992 1351 3996
rect 992 3359 1013 3363
rect 1008 3070 1012 3359
rect 1016 3077 1020 3992
rect 1345 3991 1351 3992
rect 1646 3988 1650 4009
rect 1044 3984 1637 3988
rect 1016 3073 1028 3077
rect 1008 3066 1021 3070
rect 992 3059 1014 3063
rect 1010 2770 1014 3059
rect 1017 2777 1021 3066
rect 1024 2784 1028 3073
rect 1024 2780 1032 2784
rect 1017 2773 1025 2777
rect 1010 2766 1018 2770
rect 993 2759 1011 2763
rect 1007 2471 1011 2759
rect 1014 2478 1018 2766
rect 1021 2485 1025 2773
rect 1028 2498 1032 2780
rect 1035 2498 1039 2502
rect 1028 2494 1039 2498
rect 1021 2481 1032 2485
rect 1014 2474 1025 2478
rect 1007 2467 1018 2471
rect 992 2459 1006 2463
rect 1014 2456 1018 2467
rect 1006 2452 1018 2456
rect 1006 2170 1010 2452
rect 1006 2166 1016 2170
rect 992 2159 1005 2163
rect 1012 2156 1016 2166
rect 1006 2152 1016 2156
rect 1006 1871 1010 2152
rect 1021 1925 1025 2474
rect 1028 2035 1032 2481
rect 1035 2476 1039 2494
rect 1044 2454 1048 3984
rect 1052 3956 1630 3960
rect 1052 2664 1056 3956
rect 1060 3946 1620 3949
rect 1060 3281 1063 3946
rect 1617 3935 1620 3946
rect 1626 3947 1630 3956
rect 1633 3954 1637 3984
rect 1946 3981 1950 4012
rect 2246 3974 2250 4013
rect 2546 3967 2550 4010
rect 2846 3961 2850 4013
rect 3147 3954 3151 4013
rect 1633 3950 3153 3954
rect 3447 3947 3451 4013
rect 3746 3992 3749 4012
rect 3746 3989 3752 3992
rect 1626 3943 3451 3947
rect 3749 3935 3752 3989
rect 1617 3932 3752 3935
rect 3961 3850 3965 3962
rect 1060 3278 1494 3281
rect 1491 3253 1494 3278
rect 3961 3271 3965 3846
rect 2933 3235 2990 3238
rect 2933 3230 2935 3235
rect 2940 3230 2965 3235
rect 2970 3230 2990 3235
rect 2933 3228 2990 3230
rect 3961 3134 3965 3267
rect 2920 3030 2935 3032
rect 2929 3021 2935 3030
rect 2920 2992 2935 3021
rect 3961 3003 3965 3130
rect 3961 2873 3965 2999
rect 3961 2743 3965 2869
rect 1195 2490 1199 2556
rect 1175 2459 1176 2463
rect 1039 2450 1048 2454
rect 1039 2366 1043 2450
rect 1172 2388 1176 2459
rect 1171 2376 1175 2388
rect 1028 2030 1030 2035
rect 1028 2027 1032 2030
rect 1028 2023 1034 2027
rect 1147 2024 1151 2025
rect 1021 1920 1022 1925
rect 1021 1879 1025 1920
rect 1021 1875 1027 1879
rect 1006 1867 1019 1871
rect 993 1859 1007 1863
rect 1015 1815 1019 1867
rect 1015 1807 1019 1810
rect 992 1346 1005 1350
rect 1147 1086 1151 2020
rect 1147 1052 1151 1082
rect 1154 1914 1158 1915
rect 1154 1077 1158 1910
rect 1154 1052 1158 1073
rect 1161 1804 1165 1805
rect 1161 1800 1162 1804
rect 1161 1068 1165 1800
rect 1172 1705 1176 2376
rect 1182 1904 1186 2361
rect 1172 1699 1176 1700
rect 1161 1052 1165 1064
rect 1168 1694 1172 1695
rect 1168 1059 1172 1690
rect 1195 1595 1199 2159
rect 1203 2015 1207 2659
rect 3961 2484 3965 2739
rect 3961 2375 3965 2480
rect 3961 2264 3965 2371
rect 3961 2155 3965 2260
rect 3961 2044 3965 2151
rect 3961 1934 3965 2040
rect 1168 1052 1172 1055
rect 1175 1584 1179 1585
rect 992 1046 1011 1050
rect 1175 1037 1179 1580
rect 1203 1485 1207 1859
rect 3961 1824 3965 1930
rect 3961 1715 3965 1820
rect 3961 1604 3965 1711
rect 3961 1494 3965 1600
rect 1175 1004 1179 1033
rect 1182 1474 1186 1475
rect 1182 1028 1186 1470
rect 3961 1384 3965 1490
rect 1182 1004 1186 1024
rect 1189 1364 1193 1365
rect 1189 1360 1190 1364
rect 1189 1019 1193 1360
rect 3961 1274 3965 1380
rect 1189 1004 1193 1015
rect 1196 1254 1200 1255
rect 1196 1010 1200 1250
rect 1203 1050 1207 1259
rect 3961 1150 3965 1270
rect 3968 3550 3975 3551
rect 3972 3546 3975 3550
rect 3968 3544 3975 3546
rect 3968 3235 3972 3544
rect 3968 3043 3972 3231
rect 3968 2913 3972 3039
rect 3968 2783 3972 2909
rect 3968 2654 3972 2779
rect 3968 2394 3972 2650
rect 3968 2284 3972 2390
rect 3968 2174 3972 2280
rect 3968 2064 3972 2170
rect 3968 1954 3972 2060
rect 3968 1844 3972 1950
rect 3968 1734 3972 1840
rect 3968 1624 3972 1730
rect 3968 1514 3972 1620
rect 3968 1404 3972 1510
rect 3968 1294 3972 1400
rect 3968 1184 3972 1290
rect 3968 1150 3972 1180
rect 3350 1086 3354 1087
rect 3050 1077 3054 1078
rect 2750 1068 2754 1069
rect 1203 1045 1207 1046
rect 2450 1059 2454 1060
rect 2150 1037 2154 1038
rect 1850 1028 1854 1029
rect 1550 1019 1554 1020
rect 1196 1004 1200 1006
rect 1250 1010 1254 1011
rect 1250 998 1254 1006
rect 1550 998 1554 1015
rect 1850 1000 1854 1024
rect 2150 1000 2154 1033
rect 2450 999 2454 1055
rect 2750 999 2754 1064
rect 3050 1000 3054 1073
rect 3350 1000 3354 1082
<< m3contact >>
rect 1257 4000 1266 4009
rect 1016 3992 1021 3997
rect 991 3957 1000 3966
rect 991 3657 1000 3666
rect 1006 2459 1011 2464
rect 1005 2159 1009 2163
rect 1035 2471 1040 2476
rect 1069 2985 1073 2989
rect 1231 2985 1236 2990
rect 1052 2660 1056 2664
rect 1203 2659 1208 2664
rect 1187 2487 1191 2491
rect 1170 2459 1175 2464
rect 1039 2361 1044 2366
rect 1030 2030 1035 2035
rect 1147 2020 1151 2024
rect 1022 1920 1027 1925
rect 1007 1859 1012 1864
rect 1015 1810 1020 1815
rect 1005 1346 1010 1351
rect 1036 1239 1042 1245
rect 1147 1082 1151 1086
rect 1154 1910 1158 1914
rect 1154 1073 1158 1077
rect 1162 1800 1166 1804
rect 1182 2361 1187 2366
rect 1195 2159 1200 2164
rect 1172 1700 1177 1705
rect 1161 1064 1165 1068
rect 1168 1690 1172 1694
rect 1203 2010 1208 2015
rect 1209 1900 1213 1904
rect 1203 1859 1208 1864
rect 1195 1590 1200 1595
rect 1168 1055 1172 1059
rect 1175 1580 1179 1584
rect 1211 1790 1215 1794
rect 1211 1680 1215 1684
rect 1213 1570 1217 1574
rect 1203 1480 1208 1485
rect 1175 1033 1179 1037
rect 1182 1470 1186 1474
rect 1203 1460 1207 1464
rect 1182 1024 1186 1028
rect 1190 1360 1194 1364
rect 1204 1350 1208 1354
rect 1203 1259 1208 1264
rect 1189 1015 1193 1019
rect 1196 1250 1200 1254
rect 3350 1082 3354 1086
rect 3050 1073 3054 1077
rect 2750 1064 2754 1068
rect 1203 1046 1207 1050
rect 2450 1055 2454 1059
rect 2150 1033 2154 1037
rect 1850 1024 1854 1028
rect 1550 1015 1554 1019
rect 1196 1006 1200 1010
rect 1250 1006 1254 1010
<< metal3 >>
rect 1256 4009 1267 4010
rect 1256 4007 1257 4009
rect 1046 4001 1257 4007
rect 1015 3997 1022 3998
rect 1046 3997 1052 4001
rect 1256 4000 1257 4001
rect 1266 4000 1267 4009
rect 1256 3999 1267 4000
rect 1015 3992 1016 3997
rect 1021 3992 1052 3997
rect 1015 3991 1052 3992
rect 990 3966 1001 3967
rect 990 3957 991 3966
rect 1000 3964 1001 3966
rect 1000 3958 1021 3964
rect 1000 3957 1001 3958
rect 990 3956 1001 3957
rect 990 3666 1001 3667
rect 990 3657 991 3666
rect 1000 3664 1001 3666
rect 1000 3658 1012 3664
rect 1000 3657 1001 3658
rect 990 3656 1001 3657
rect 1006 2492 1012 3658
rect 1015 2557 1021 3958
rect 3655 3549 3738 3557
rect 3641 3542 3738 3549
rect 3641 3535 3748 3542
rect 3804 3541 3848 3552
rect 3624 3533 3748 3535
rect 3624 3525 3679 3533
rect 3618 3511 3665 3525
rect 3714 3519 3748 3533
rect 3773 3526 3848 3541
rect 3773 3525 3865 3526
rect 3754 3519 3865 3525
rect 3714 3518 3865 3519
rect 3724 3517 3865 3518
rect 3618 3501 3648 3511
rect 3724 3501 3797 3517
rect 3824 3502 3865 3517
rect 3618 3466 3642 3501
rect 3724 3495 3778 3501
rect 3731 3492 3778 3495
rect 3841 3487 3865 3502
rect 3618 3455 3653 3466
rect 3618 3442 3658 3455
rect 3629 3441 3658 3442
rect 3841 3444 3871 3487
rect 3629 3431 3668 3441
rect 3841 3440 3865 3444
rect 3634 3429 3668 3431
rect 3634 3417 3679 3429
rect 3830 3428 3865 3440
rect 3644 3414 3679 3417
rect 3824 3416 3865 3428
rect 3824 3415 3854 3416
rect 3644 3406 3690 3414
rect 3644 3405 3697 3406
rect 3655 3403 3697 3405
rect 3798 3404 3854 3415
rect 3655 3390 3700 3403
rect 3798 3400 3848 3404
rect 3666 3381 3700 3390
rect 3765 3391 3848 3400
rect 3765 3387 3822 3391
rect 3670 3360 3703 3381
rect 3750 3376 3822 3387
rect 3750 3370 3789 3376
rect 3732 3363 3789 3370
rect 3670 3358 3726 3360
rect 3732 3358 3774 3363
rect 3670 3357 3774 3358
rect 3679 3346 3774 3357
rect 3679 3336 3756 3346
rect 3691 3334 3756 3336
rect 3691 3327 3736 3334
rect 3689 3305 3736 3327
rect 3689 3293 3725 3305
rect 1230 2990 1237 2991
rect 1068 2989 1231 2990
rect 1068 2985 1069 2989
rect 1073 2985 1231 2989
rect 1236 2985 1237 2990
rect 1068 2984 1237 2985
rect 1051 2664 1209 2665
rect 1051 2660 1052 2664
rect 1056 2660 1203 2664
rect 1051 2659 1203 2660
rect 1208 2659 1209 2664
rect 1202 2658 1209 2659
rect 1015 2551 1200 2557
rect 1006 2491 1192 2492
rect 1006 2487 1187 2491
rect 1191 2487 1192 2491
rect 1006 2486 1192 2487
rect 1034 2476 1041 2477
rect 1034 2471 1035 2476
rect 1040 2471 1184 2476
rect 1034 2470 1184 2471
rect 1005 2464 1012 2465
rect 1169 2464 1176 2465
rect 1005 2459 1006 2464
rect 1011 2459 1170 2464
rect 1175 2459 1178 2464
rect 1005 2458 1178 2459
rect 1178 2379 1179 2380
rect 1038 2366 1045 2367
rect 1181 2366 1188 2367
rect 1038 2361 1039 2366
rect 1044 2361 1182 2366
rect 1187 2361 1188 2366
rect 1038 2360 1188 2361
rect 1194 2164 1201 2165
rect 1004 2163 1195 2164
rect 1004 2159 1005 2163
rect 1009 2159 1195 2163
rect 1200 2159 1212 2164
rect 1004 2158 1212 2159
rect 1029 2035 1036 2036
rect 1027 2030 1030 2035
rect 1035 2030 1202 2035
rect 1027 2029 1202 2030
rect 1146 2024 1206 2025
rect 1146 2020 1147 2024
rect 1151 2020 1206 2024
rect 1146 2019 1206 2020
rect 1202 2015 1209 2016
rect 1202 2010 1203 2015
rect 1208 2010 1209 2015
rect 1202 2009 1209 2010
rect 1021 1925 1028 1926
rect 1021 1920 1022 1925
rect 1027 1920 1202 1925
rect 1021 1919 1202 1920
rect 1153 1914 1204 1915
rect 1153 1910 1154 1914
rect 1158 1910 1204 1914
rect 1153 1909 1204 1910
rect 1006 1864 1013 1865
rect 1202 1864 1209 1865
rect 1006 1859 1007 1864
rect 1012 1859 1203 1864
rect 1208 1859 1212 1864
rect 1006 1858 1212 1859
rect 1014 1815 1021 1816
rect 1014 1810 1015 1815
rect 1020 1810 1202 1815
rect 1014 1809 1202 1810
rect 1161 1804 1207 1805
rect 1161 1800 1162 1804
rect 1166 1800 1207 1804
rect 1161 1799 1207 1800
rect 1171 1705 1178 1706
rect 1171 1700 1172 1705
rect 1177 1700 1202 1705
rect 1171 1699 1202 1700
rect 1167 1694 1203 1695
rect 1167 1690 1168 1694
rect 1172 1690 1203 1694
rect 1167 1689 1203 1690
rect 1194 1595 1201 1596
rect 1194 1590 1195 1595
rect 1200 1590 1202 1595
rect 1194 1589 1202 1590
rect 1174 1584 1202 1585
rect 1174 1580 1175 1584
rect 1179 1580 1202 1584
rect 1174 1579 1202 1580
rect 1202 1485 1209 1486
rect 1202 1480 1203 1485
rect 1208 1480 1209 1485
rect 1202 1479 1209 1480
rect 1181 1474 1202 1475
rect 1181 1470 1182 1474
rect 1186 1470 1202 1474
rect 1181 1469 1202 1470
rect 1181 1369 1206 1375
rect 1181 1365 1186 1369
rect 1132 1359 1186 1365
rect 1189 1364 1203 1365
rect 1189 1360 1190 1364
rect 1194 1360 1203 1364
rect 1189 1359 1203 1360
rect 1004 1351 1011 1352
rect 1132 1351 1138 1359
rect 1004 1346 1005 1351
rect 1010 1346 1138 1351
rect 1004 1345 1138 1346
rect 1202 1264 1209 1265
rect 1202 1259 1203 1264
rect 1208 1259 1209 1264
rect 1202 1258 1209 1259
rect 1194 1254 1205 1255
rect 1194 1250 1196 1254
rect 1200 1250 1205 1254
rect 1194 1249 1205 1250
rect 1035 1245 1043 1246
rect 1035 1239 1036 1245
rect 1042 1239 1206 1245
rect 1035 1238 1043 1239
rect 1144 1086 3362 1087
rect 1144 1082 1147 1086
rect 1151 1082 3350 1086
rect 3354 1082 3362 1086
rect 1144 1081 3362 1082
rect 1144 1077 3065 1078
rect 1144 1073 1154 1077
rect 1158 1073 3050 1077
rect 3054 1073 3065 1077
rect 1144 1072 3065 1073
rect 1144 1068 2760 1069
rect 1144 1064 1161 1068
rect 1165 1064 2750 1068
rect 2754 1064 2760 1068
rect 1144 1063 2760 1064
rect 1144 1059 2465 1060
rect 1144 1055 1168 1059
rect 1172 1055 2450 1059
rect 2454 1055 2465 1059
rect 1144 1054 2465 1055
rect 1005 1050 1211 1051
rect 1005 1046 1203 1050
rect 1207 1046 1211 1050
rect 1005 1045 1211 1046
rect 1153 1037 2165 1038
rect 1153 1033 1175 1037
rect 1179 1033 2150 1037
rect 2154 1033 2165 1037
rect 1153 1032 2165 1033
rect 1153 1028 1859 1029
rect 1153 1024 1182 1028
rect 1186 1024 1850 1028
rect 1854 1024 1859 1028
rect 1153 1023 1859 1024
rect 1153 1019 1560 1020
rect 1153 1015 1189 1019
rect 1193 1015 1550 1019
rect 1554 1015 1560 1019
rect 1153 1014 1560 1015
rect 1153 1010 1351 1011
rect 1153 1006 1196 1010
rect 1200 1006 1250 1010
rect 1254 1006 1351 1010
rect 1153 1005 1351 1006
<< m2p >>
rect 1002 1859 1003 1863
use PADFC  PADFC_0
timestamp 949001400
transform 1 0 0 0 1 4000
box 327 -3 1003 673
use PADINC  reset
timestamp 1084294328
transform 1 0 1000 0 1 4000
box -6 -3 303 1000
use PADOUT  adr0
timestamp 1084294529
transform 1 0 1300 0 1 4000
box -6 -3 303 1000
use PADOUT  adr1
timestamp 1084294529
transform 1 0 1600 0 1 4000
box -6 -3 303 1000
use PADOUT  adr2
timestamp 1084294529
transform 1 0 1900 0 1 4000
box -6 -3 303 1000
use PADOUT  adr3
timestamp 1084294529
transform 1 0 2200 0 1 4000
box -6 -3 303 1000
use PADOUT  adr4
timestamp 1084294529
transform 1 0 2500 0 1 4000
box -6 -3 303 1000
use PADOUT  adr5
timestamp 1084294529
transform 1 0 2800 0 1 4000
box -6 -3 303 1000
use PADOUT  adr6
timestamp 1084294529
transform 1 0 3100 0 1 4000
box -6 -3 303 1000
use PADOUT  adr7
timestamp 1084294529
transform 1 0 3400 0 1 4000
box -6 -3 303 1000
use PADOUT  MemWrite
timestamp 1084294529
transform 1 0 3700 0 1 4000
box -6 -3 303 1000
use PADFC  PADFC_3
timestamp 949001400
transform 0 1 4000 -1 0 5000
box 327 -3 1003 673
use PADINC  ph1
timestamp 1084294328
transform 0 -1 1000 1 0 3700
box -6 -3 303 1000
use PADINC  ph2
timestamp 1084294328
transform 0 -1 1000 1 0 3400
box -6 -3 303 1000
use PADVDD  PADVDD_0
timestamp 1084294447
transform 0 1 4000 -1 0 3997
box -3 -3 303 1000
use PADGND  PADGND_0
timestamp 1084294269
transform 0 1 4000 -1 0 3698
box -3 -3 303 1000
use PADINC  memdata7
timestamp 1084294328
transform 0 -1 1000 1 0 3100
box -6 -3 303 1000
use PADINC  memdata6
timestamp 1084294328
transform 0 -1 1000 1 0 2800
box -6 -3 303 1000
use PADINC  memdata5
timestamp 1084294328
transform 0 -1 1000 1 0 2500
box -6 -3 303 1000
use PADINC  memdata4
timestamp 1084294328
transform 0 -1 1000 1 0 2200
box -6 -3 303 1000
use PADINC  memdata3
timestamp 1084294328
transform 0 -1 1000 1 0 1900
box -6 -3 303 1000
use PADINC  memdata2
timestamp 1084294328
transform 0 -1 1000 1 0 1600
box -6 -3 303 1000
use PADOUT  memdata1
timestamp 1084294529
transform 0 -1 1000 1 0 1300
box -6 -3 303 1000
use datapath  datapath_0
timestamp 1494282038
transform 1 0 1219 0 1 1182
box -168 -32 2739 2085
use PADNC  PADNC_9
timestamp 1084294400
transform 0 1 4000 1 0 3100
box -3 -3 303 1000
use PADNC  PADNC_8
timestamp 1084294400
transform 0 1 4000 1 0 2800
box -3 -3 303 1000
use PADNC  PADNC_7
timestamp 1084294400
transform 0 1 4000 1 0 2500
box -3 -3 303 1000
use PADNC  PADNC_6
timestamp 1084294400
transform 0 1 4000 1 0 2200
box -3 -3 303 1000
use PADNC  PADNC_5
timestamp 1084294400
transform 0 1 4000 1 0 1900
box -3 -3 303 1000
use PADNC  PADNC_4
timestamp 1084294400
transform 0 1 4000 1 0 1600
box -3 -3 303 1000
use PADNC  PADNC_3
timestamp 1084294400
transform 0 1 4000 1 0 1300
box -3 -3 303 1000
use PADOUT  memdata0
timestamp 1084294529
transform 0 -1 1000 1 0 1000
box -6 -3 303 1000
use PADFC  PADFC_2
timestamp 949001400
transform 0 -1 1000 1 0 0
box 327 -3 1003 673
use PADOUT  writedata0
timestamp 1084294529
transform -1 0 1300 0 -1 1000
box -6 -3 303 1000
use PADOUT  writedata1
timestamp 1084294529
transform -1 0 1600 0 -1 1000
box -6 -3 303 1000
use PADOUT  writedata2
timestamp 1084294529
transform -1 0 1900 0 -1 1000
box -6 -3 303 1000
use PADOUT  writedata3
timestamp 1084294529
transform -1 0 2200 0 -1 1000
box -6 -3 303 1000
use PADOUT  writedata4
timestamp 1084294529
transform -1 0 2500 0 -1 1000
box -6 -3 303 1000
use PADOUT  writedata5
timestamp 1084294529
transform -1 0 2800 0 -1 1000
box -6 -3 303 1000
use PADOUT  writedata6
timestamp 1084294529
transform -1 0 3100 0 -1 1000
box -6 -3 303 1000
use PADOUT  writedata7
timestamp 1084294529
transform -1 0 3400 0 -1 1000
box -6 -3 303 1000
use PADNC  PADNC_0
timestamp 1084294400
transform 1 0 3400 0 -1 1000
box -3 -3 303 1000
use PADNC  PADNC_1
timestamp 1084294400
transform 0 1 4000 1 0 1000
box -3 -3 303 1000
use PADFC  PADFC_1
timestamp 949001400
transform -1 0 4998 0 -1 1000
box 327 -3 1003 673
use PADNC  PADNC_2
timestamp 1084294400
transform 1 0 3700 0 -1 1000
box -3 -3 303 1000
<< end >>
