magic
tech scmos
timestamp 1490727624
<< m2contact >>
rect -2 -2 2 2
<< end >>
