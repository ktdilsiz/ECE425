magic
tech scmos
timestamp 1487715963
<< nwell >>
rect -6 40 50 96
<< ntransistor >>
rect 5 26 7 30
rect 10 26 12 30
rect 18 26 20 30
rect 23 26 25 30
rect 31 26 33 30
<< ptransistor >>
rect 35 76 39 78
rect 5 54 7 58
rect 13 54 15 58
rect 21 54 23 58
rect 29 54 31 58
<< ndiffusion >>
rect 4 26 5 30
rect 7 26 10 30
rect 12 26 13 30
rect 17 26 18 30
rect 20 26 23 30
rect 25 26 26 30
rect 30 26 31 30
rect 33 26 34 30
<< pdiffusion >>
rect 35 78 39 79
rect 35 75 39 76
rect 4 54 5 58
rect 7 54 8 58
rect 12 54 13 58
rect 15 54 16 58
rect 20 54 21 58
rect 23 54 24 58
rect 28 54 29 58
rect 31 54 32 58
<< ndcontact >>
rect 0 26 4 30
rect 13 26 17 30
rect 26 26 30 30
rect 34 26 38 30
<< pdcontact >>
rect 35 79 39 83
rect 35 71 39 75
rect 0 54 4 58
rect 8 54 12 58
rect 16 54 20 58
rect 24 54 28 58
rect 32 54 36 58
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
rect 40 -2 44 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
rect 32 88 36 92
rect 40 88 44 92
<< polysilicon >>
rect 33 76 35 78
rect 39 76 42 78
rect 5 58 7 60
rect 13 58 15 60
rect 21 58 23 60
rect 29 58 31 60
rect 5 53 7 54
rect 13 53 15 54
rect 21 53 23 54
rect 2 51 7 53
rect 10 51 15 53
rect 18 51 23 53
rect 29 53 31 54
rect 29 51 34 53
rect 2 44 4 51
rect 10 44 12 51
rect 18 44 20 51
rect 32 48 34 51
rect 2 33 4 40
rect 2 31 7 33
rect 5 30 7 31
rect 10 30 12 40
rect 18 30 20 40
rect 26 45 32 47
rect 26 35 28 45
rect 23 33 28 35
rect 31 33 32 35
rect 40 36 42 76
rect 36 34 42 36
rect 23 30 25 33
rect 31 30 33 33
rect 5 24 7 26
rect 10 24 12 26
rect 18 24 20 26
rect 23 24 25 26
rect 31 24 33 26
<< polycontact >>
rect 0 40 4 44
rect 8 40 12 44
rect 16 40 20 44
rect 32 44 36 48
rect 32 33 36 37
<< metal1 >>
rect -2 92 46 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 32 92
rect 36 88 40 92
rect 44 88 46 92
rect -2 86 46 88
rect 8 58 12 86
rect 35 83 39 86
rect 35 78 39 79
rect 39 71 44 75
rect 16 61 36 65
rect 16 58 20 61
rect 32 58 36 61
rect 0 51 4 54
rect 16 51 20 54
rect 0 47 20 51
rect 24 37 28 54
rect 40 44 44 71
rect 13 33 32 37
rect 13 30 17 33
rect 40 30 44 40
rect 38 26 44 30
rect 0 4 4 26
rect 26 4 30 26
rect -2 2 46 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 40 2
rect 44 -2 46 2
rect -2 -4 46 -2
<< m2contact >>
rect 0 40 4 44
rect 8 40 12 44
rect 16 40 20 44
rect 32 44 36 48
rect 40 40 44 44
<< labels >>
rlabel metal1 -1 0 -1 0 2 Gnd!
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel m2contact 2 42 2 42 1 a
rlabel m2contact 10 42 10 42 1 b
rlabel m2contact 18 42 18 42 1 c
rlabel m2contact 34 46 34 46 1 d
rlabel m2contact 42 42 42 42 1 y
<< end >>
