magic
tech scmos
timestamp 1488311641
<< m2contact >>
rect -2 -2 2 2
<< end >>
