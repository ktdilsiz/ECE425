magic
tech scmos
timestamp 1484533408
<< nwell >>
rect -6 40 50 96
<< ntransistor >>
rect 5 7 7 31
rect 10 7 12 31
rect 15 7 17 31
rect 20 7 22 31
rect 25 7 27 31
<< ptransistor >>
rect 5 68 7 83
rect 13 68 15 83
rect 21 68 23 83
rect 29 68 31 83
rect 37 68 39 83
<< ndiffusion >>
rect 4 7 5 31
rect 7 7 10 31
rect 12 7 15 31
rect 17 7 20 31
rect 22 7 25 31
rect 27 7 28 31
<< pdiffusion >>
rect 0 82 5 83
rect 4 68 5 82
rect 7 82 13 83
rect 7 68 8 82
rect 12 68 13 82
rect 15 82 21 83
rect 15 68 16 82
rect 20 68 21 82
rect 23 82 29 83
rect 23 68 24 82
rect 28 68 29 82
rect 31 82 37 83
rect 31 68 32 82
rect 36 68 37 82
rect 39 82 44 83
rect 39 68 40 82
<< ndcontact >>
rect 0 7 4 31
rect 28 7 32 31
<< pdcontact >>
rect 0 68 4 82
rect 8 68 12 82
rect 16 68 20 82
rect 24 68 28 82
rect 32 68 36 82
rect 40 68 44 82
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
rect 40 -2 44 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
rect 32 88 36 92
rect 40 88 44 92
<< polysilicon >>
rect 5 83 7 85
rect 13 83 15 85
rect 21 83 23 85
rect 29 83 31 85
rect 37 83 39 85
rect 5 60 7 68
rect 13 67 15 68
rect 0 58 7 60
rect 10 65 15 67
rect 0 57 4 58
rect 0 39 2 53
rect 0 37 7 39
rect 5 31 7 37
rect 10 31 12 65
rect 21 48 23 68
rect 15 44 16 48
rect 20 46 23 48
rect 15 31 17 44
rect 29 40 31 68
rect 37 60 39 68
rect 37 58 44 60
rect 40 57 44 58
rect 20 38 31 40
rect 20 31 22 38
rect 42 35 44 53
rect 25 33 44 35
rect 25 31 27 33
rect 5 5 7 7
rect 10 5 12 7
rect 15 5 17 7
rect 20 5 22 7
rect 25 5 27 7
<< polycontact >>
rect 0 53 4 57
rect 6 44 10 48
rect 16 44 20 48
rect 40 53 44 57
rect 31 44 35 48
<< metal1 >>
rect -2 92 46 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 32 92
rect 36 88 40 92
rect 44 88 46 92
rect -2 86 46 88
rect 0 82 4 86
rect 8 82 12 83
rect 16 82 20 86
rect 24 82 28 83
rect 32 82 36 86
rect 40 82 44 83
rect 8 57 12 68
rect 24 64 28 68
rect 40 64 44 68
rect 24 60 44 64
rect 24 57 28 60
rect 8 53 24 57
rect 24 39 28 53
rect 24 35 32 39
rect 28 31 32 35
rect 0 4 4 7
rect -2 2 46 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 40 2
rect 44 -2 46 2
rect -2 -4 46 -2
<< m2contact >>
rect 0 53 4 57
rect 24 53 28 57
rect 40 53 44 57
rect 8 44 10 48
rect 10 44 12 48
rect 16 44 20 48
rect 32 44 35 48
rect 35 44 36 48
<< labels >>
rlabel metal1 -1 0 -1 0 2 Gnd!
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel m2contact 2 55 2 55 1 a
rlabel m2contact 10 46 10 46 1 b
rlabel m2contact 18 46 18 46 1 c
rlabel m2contact 26 55 26 55 1 y
rlabel m2contact 42 55 42 55 1 e
rlabel m2contact 34 46 34 46 1 d
<< end >>
