magic
tech scmos
timestamp 1488311641
<< m2contact >>
rect -7 -7 7 7
<< end >>
