magic
tech scmos
timestamp 1489950195
<< nwell >>
rect -6 40 34 96
<< ntransistor >>
rect 5 7 7 21
rect 13 7 15 21
rect 21 7 23 21
<< ptransistor >>
rect 5 63 7 83
rect 10 63 12 83
rect 18 73 20 83
<< ndiffusion >>
rect 4 7 5 21
rect 7 7 8 21
rect 12 7 13 21
rect 15 7 16 21
rect 20 7 21 21
rect 23 7 24 21
<< pdiffusion >>
rect 0 82 5 83
rect 4 63 5 82
rect 7 63 10 83
rect 12 82 18 83
rect 12 63 13 82
rect 17 73 18 82
rect 20 82 25 83
rect 20 73 21 82
<< ndcontact >>
rect 0 7 4 21
rect 8 7 12 21
rect 16 7 20 21
rect 24 7 28 21
<< pdcontact >>
rect 0 63 4 82
rect 13 63 17 82
rect 21 73 25 82
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
<< polysilicon >>
rect 5 83 7 85
rect 10 83 12 85
rect 18 83 20 85
rect 5 62 7 63
rect 1 60 7 62
rect 1 45 3 60
rect 10 45 12 63
rect 1 24 3 41
rect 10 24 12 41
rect 18 24 20 73
rect 1 22 7 24
rect 10 22 15 24
rect 18 22 23 24
rect 5 21 7 22
rect 13 21 15 22
rect 21 21 23 22
rect 5 5 7 7
rect 13 5 15 7
rect 21 5 23 7
<< polycontact >>
rect 0 41 4 45
rect 9 41 13 45
rect 20 58 24 62
<< metal1 >>
rect -2 92 30 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 30 92
rect -2 86 30 88
rect 0 82 4 86
rect 13 82 17 83
rect 21 82 25 86
rect 13 52 17 63
rect 13 48 16 52
rect 20 48 28 52
rect 0 25 20 29
rect 0 21 4 25
rect 16 21 20 25
rect 24 21 28 48
rect 8 4 12 7
rect -2 2 30 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 30 2
rect -2 -4 30 -2
<< m2contact >>
rect 24 58 28 62
rect 16 48 20 52
rect 0 41 4 45
rect 8 41 9 45
rect 9 41 12 45
<< labels >>
rlabel m2contact 2 43 2 43 1 a
rlabel m2contact 10 43 10 43 1 b
rlabel m2contact 18 50 18 50 1 y
rlabel m2contact 26 60 26 60 1 c
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel metal1 -1 0 -1 0 2 Gnd!
<< end >>
