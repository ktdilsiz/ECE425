magic
tech scmos
timestamp 1493754926
<< metal1 >>
rect 6 966 62 974
rect 20 918 27 922
rect 6 876 62 884
rect 52 868 56 872
rect 84 868 88 872
rect 116 868 120 872
<< m2contact >>
rect 16 918 20 922
rect 32 918 36 922
rect 48 918 52 922
rect 48 868 52 872
rect 56 868 60 872
rect 80 868 84 872
rect 88 868 92 872
rect 112 868 116 872
rect 120 868 124 872
<< metal2 >>
rect -1 932 5 933
rect -1 928 0 932
rect 4 928 5 932
rect -1 927 5 928
rect 15 932 21 933
rect 15 928 16 932
rect 20 928 21 932
rect 15 927 21 928
rect 0 63 4 927
rect 16 922 20 927
rect 32 913 36 918
rect 7 912 13 913
rect 7 908 8 912
rect 12 908 13 912
rect 7 907 13 908
rect 31 912 37 913
rect 31 908 32 912
rect 36 908 37 912
rect 31 907 37 908
rect 8 36 12 907
rect 48 893 52 918
rect 103 912 109 913
rect 103 908 104 912
rect 108 908 109 912
rect 103 907 109 908
rect 135 912 141 913
rect 135 908 136 912
rect 140 908 141 912
rect 135 907 141 908
rect 15 892 21 893
rect 15 888 16 892
rect 20 888 21 892
rect 15 887 21 888
rect 47 892 53 893
rect 47 888 48 892
rect 52 888 53 892
rect 47 887 53 888
rect 16 54 20 887
rect 56 872 60 878
rect 88 872 92 878
rect 48 44 52 868
rect 80 54 84 868
rect 104 26 108 907
rect 120 872 124 878
rect 136 874 140 907
rect 112 54 116 868
<< m3contact >>
rect 0 928 4 932
rect 16 928 20 932
rect 8 908 12 912
rect 32 908 36 912
rect 104 908 108 912
rect 136 908 140 912
rect 16 888 20 892
rect 48 888 52 892
<< metal3 >>
rect -1 932 21 933
rect -1 928 0 932
rect 4 928 16 932
rect 20 928 21 932
rect -1 927 21 928
rect 7 912 37 913
rect 7 908 8 912
rect 12 908 32 912
rect 36 908 37 912
rect 7 907 37 908
rect 103 912 141 913
rect 103 908 104 912
rect 108 908 136 912
rect 140 908 141 912
rect 103 907 141 908
rect 15 892 53 893
rect 15 888 16 892
rect 20 888 48 892
rect 52 888 53 892
rect 15 887 53 888
use inv_4x  inv_4x_0
timestamp 1484455226
transform 1 0 8 0 1 880
box -6 -4 18 96
use inv_4x  inv_4x_1
timestamp 1484455226
transform 1 0 24 0 1 880
box -6 -4 18 96
use inv_4x  inv_4x_2
timestamp 1484455226
transform 1 0 40 0 1 880
box -6 -4 18 96
use clkinvbufdual_4x  clkinvbufdual_4x_0
timestamp 1484532171
transform 1 0 56 0 1 880
box -6 -6 90 96
use flopenr_dp_1x  flopenr_dp_1x_0
timestamp 1493662838
transform 1 0 0 0 1 770
box -6 -4 147 96
use flopenr_dp_1x  flopenr_dp_1x_1
timestamp 1493662838
transform 1 0 0 0 1 660
box -6 -4 147 96
use flopenr_dp_1x  flopenr_dp_1x_2
timestamp 1493662838
transform 1 0 0 0 1 550
box -6 -4 147 96
use flopenr_dp_1x  flopenr_dp_1x_3
timestamp 1493662838
transform 1 0 0 0 1 440
box -6 -4 147 96
use flopenr_dp_1x  flopenr_dp_1x_4
timestamp 1493662838
transform 1 0 0 0 1 330
box -6 -4 147 96
use flopenr_dp_1x  flopenr_dp_1x_5
timestamp 1493662838
transform 1 0 0 0 1 220
box -6 -4 147 96
use flopenr_dp_1x  flopenr_dp_1x_6
timestamp 1493662838
transform 1 0 0 0 1 110
box -6 -4 147 96
use flopenr_dp_1x  flopenr_dp_1x_7
timestamp 1493662838
transform 1 0 0 0 1 0
box -6 -4 147 96
<< end >>
