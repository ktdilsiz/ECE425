magic
tech scmos
timestamp 1484455043
<< nwell >>
rect -6 40 138 96
<< ntransistor >>
rect 11 8 13 26
rect 19 8 21 14
rect 27 8 29 14
rect 32 8 34 14
rect 53 8 55 14
rect 61 8 63 12
rect 68 8 70 12
rect 77 8 79 14
rect 85 8 87 14
rect 93 8 95 12
rect 100 8 102 12
rect 109 8 111 14
rect 125 8 127 15
<< ptransistor >>
rect 5 71 7 83
rect 10 71 12 83
rect 18 77 20 83
rect 23 77 25 83
rect 53 77 55 83
rect 61 79 63 83
rect 68 79 70 83
rect 77 74 79 83
rect 85 77 87 83
rect 93 79 95 83
rect 100 79 102 83
rect 109 74 111 83
rect 125 73 127 83
<< ndiffusion >>
rect 6 24 11 26
rect 10 10 11 24
rect 6 8 11 10
rect 13 24 18 26
rect 13 10 14 24
rect 18 10 19 14
rect 13 8 19 10
rect 21 13 27 14
rect 21 9 22 13
rect 26 9 27 13
rect 21 8 27 9
rect 29 8 32 14
rect 34 13 39 14
rect 34 9 35 13
rect 34 8 39 9
rect 52 8 53 14
rect 55 8 56 14
rect 72 13 77 14
rect 60 8 61 12
rect 63 8 68 12
rect 70 9 72 12
rect 76 9 77 13
rect 70 8 77 9
rect 79 8 80 14
rect 84 8 85 14
rect 87 8 88 14
rect 104 13 109 14
rect 92 8 93 12
rect 95 8 100 12
rect 102 9 104 12
rect 108 9 109 13
rect 102 8 109 9
rect 111 8 112 14
rect 120 13 125 15
rect 124 9 125 13
rect 120 8 125 9
rect 127 13 132 15
rect 127 9 128 13
rect 127 8 132 9
<< pdiffusion >>
rect 0 81 5 83
rect 4 72 5 81
rect 0 71 5 72
rect 7 71 10 83
rect 12 81 18 83
rect 12 72 13 81
rect 17 77 18 81
rect 20 77 23 83
rect 25 82 30 83
rect 25 78 26 82
rect 25 77 30 78
rect 48 82 53 83
rect 52 78 53 82
rect 48 77 53 78
rect 55 77 56 83
rect 60 79 61 83
rect 63 79 68 83
rect 70 79 72 83
rect 12 71 17 72
rect 76 74 77 83
rect 79 74 80 83
rect 84 77 85 83
rect 87 77 88 83
rect 92 79 93 83
rect 95 79 100 83
rect 102 79 104 83
rect 108 74 109 83
rect 111 74 112 83
rect 120 82 125 83
rect 124 73 125 82
rect 127 82 132 83
rect 127 73 128 82
<< ndcontact >>
rect 6 10 10 24
rect 14 10 18 24
rect 22 9 26 13
rect 35 9 39 13
rect 48 8 52 14
rect 56 8 60 14
rect 72 9 76 13
rect 80 8 84 14
rect 88 8 92 14
rect 104 9 108 13
rect 112 8 116 14
rect 120 9 124 13
rect 128 9 132 13
<< pdcontact >>
rect 0 72 4 81
rect 13 72 17 81
rect 26 78 30 82
rect 48 78 52 82
rect 56 77 60 83
rect 72 74 76 83
rect 80 74 84 83
rect 88 77 92 83
rect 104 74 108 83
rect 112 74 116 83
rect 120 73 124 82
rect 128 73 132 82
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
rect 40 -2 44 2
rect 48 -2 52 2
rect 56 -2 60 2
rect 64 -2 68 2
rect 72 -2 76 2
rect 80 -2 84 2
rect 88 -2 92 2
rect 96 -2 100 2
rect 104 -2 108 2
rect 112 -2 116 2
rect 120 -2 124 2
rect 128 -2 132 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
rect 32 88 36 92
rect 40 88 44 92
rect 48 88 52 92
rect 56 88 60 92
rect 64 88 68 92
rect 72 88 76 92
rect 80 88 84 92
rect 88 88 92 92
rect 96 88 100 92
rect 104 88 108 92
rect 112 88 116 92
rect 120 88 124 92
rect 128 88 132 92
<< polysilicon >>
rect 5 83 7 85
rect 10 83 12 85
rect 18 83 20 85
rect 23 83 25 85
rect 53 83 55 85
rect 61 83 63 85
rect 68 83 70 85
rect 77 83 79 85
rect 85 83 87 85
rect 93 83 95 85
rect 100 83 102 85
rect 109 83 111 85
rect 125 83 127 85
rect 5 66 7 71
rect 4 64 7 66
rect 10 66 12 71
rect 10 64 15 66
rect 13 47 15 64
rect 18 55 20 77
rect 23 61 25 77
rect 23 59 31 61
rect 18 53 26 55
rect 16 43 21 46
rect 11 26 13 35
rect 19 14 21 43
rect 24 36 26 53
rect 29 49 31 59
rect 53 57 55 77
rect 61 74 63 79
rect 68 67 70 79
rect 68 63 69 67
rect 29 47 32 49
rect 53 45 55 53
rect 53 43 63 45
rect 24 34 48 36
rect 27 14 29 34
rect 32 26 33 29
rect 32 14 34 26
rect 53 14 55 17
rect 61 12 63 43
rect 68 12 70 63
rect 77 28 79 74
rect 85 57 87 77
rect 93 74 95 79
rect 100 67 102 79
rect 100 63 101 67
rect 88 53 95 55
rect 78 24 79 28
rect 77 14 79 24
rect 85 14 87 17
rect 93 12 95 53
rect 100 12 102 63
rect 109 36 111 74
rect 110 32 111 36
rect 109 14 111 32
rect 125 15 127 73
rect 11 6 13 8
rect 19 6 21 8
rect 27 6 29 8
rect 32 6 34 8
rect 53 6 55 8
rect 61 6 63 8
rect 68 6 70 8
rect 77 6 79 8
rect 85 6 87 8
rect 93 6 95 8
rect 100 6 102 8
rect 109 6 111 8
rect 125 6 127 8
<< polycontact >>
rect 0 62 4 66
rect 12 43 16 47
rect 11 35 15 39
rect 60 70 64 74
rect 69 63 73 67
rect 52 53 56 57
rect 32 45 36 49
rect 48 33 52 37
rect 33 26 37 30
rect 52 17 56 21
rect 92 70 96 74
rect 101 63 105 67
rect 84 53 88 57
rect 74 24 78 28
rect 84 17 88 21
rect 121 39 125 43
rect 106 32 110 36
<< metal1 >>
rect -2 92 134 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 32 92
rect 36 88 40 92
rect 44 88 48 92
rect 52 88 56 92
rect 60 88 64 92
rect 68 88 72 92
rect 76 88 80 92
rect 84 88 88 92
rect 92 88 96 92
rect 100 88 104 92
rect 108 88 112 92
rect 116 88 120 92
rect 124 88 128 92
rect 132 88 134 92
rect -2 86 134 88
rect 0 81 4 86
rect 0 71 4 72
rect 13 81 17 83
rect 26 82 30 86
rect 72 83 76 86
rect 104 83 108 86
rect 26 77 30 78
rect 48 82 52 83
rect 17 72 24 74
rect 13 70 24 72
rect 28 71 37 74
rect 48 71 52 78
rect 28 70 48 71
rect 33 67 48 70
rect 80 67 84 74
rect 112 67 116 74
rect 120 82 124 86
rect 128 82 132 83
rect 4 62 32 64
rect 0 60 32 62
rect 73 63 80 67
rect 105 63 116 67
rect 56 53 72 57
rect 88 53 104 57
rect 32 39 36 45
rect 112 43 116 63
rect 128 46 132 73
rect 116 39 121 43
rect 15 35 36 39
rect 52 33 88 37
rect 92 36 93 37
rect 92 33 106 36
rect 88 32 106 33
rect 6 24 10 26
rect 6 4 10 10
rect 14 24 18 26
rect 60 24 74 28
rect 96 21 100 25
rect 14 8 18 10
rect 22 16 24 19
rect 56 17 64 21
rect 88 17 100 21
rect 22 15 28 16
rect 22 13 26 15
rect 22 8 26 9
rect 35 13 39 14
rect 35 4 39 9
rect 72 13 76 14
rect 72 4 76 9
rect 104 13 108 14
rect 104 4 108 9
rect 120 13 124 15
rect 120 4 124 9
rect 128 13 132 42
rect 128 8 132 9
rect -2 2 134 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 40 2
rect 44 -2 48 2
rect 52 -2 56 2
rect 60 -2 64 2
rect 68 -2 72 2
rect 76 -2 80 2
rect 84 -2 88 2
rect 92 -2 96 2
rect 100 -2 104 2
rect 108 -2 112 2
rect 116 -2 120 2
rect 124 -2 128 2
rect 132 -2 134 2
rect -2 -4 134 -2
<< m2contact >>
rect 24 70 28 74
rect 56 77 60 81
rect 88 77 92 81
rect 48 67 52 71
rect 64 70 68 74
rect 96 70 100 74
rect 0 62 4 66
rect 32 60 36 64
rect 80 63 84 67
rect 72 53 76 57
rect 104 53 108 57
rect 16 43 20 47
rect 64 43 68 47
rect 112 39 116 43
rect 128 42 132 46
rect 8 35 11 39
rect 11 35 12 39
rect 88 33 92 37
rect 32 26 33 30
rect 33 26 36 30
rect 56 24 60 28
rect 96 25 100 29
rect 24 16 28 20
rect 64 17 68 21
rect 48 10 52 14
rect 56 10 60 14
rect 80 10 84 14
rect 88 10 92 14
rect 112 10 116 14
<< metal2 >>
rect 24 20 28 70
rect 32 30 36 60
rect 48 14 52 67
rect 56 28 60 77
rect 56 14 60 24
rect 64 47 68 70
rect 64 21 68 43
rect 80 14 84 63
rect 88 37 92 77
rect 88 14 92 33
rect 96 29 100 70
rect 112 14 116 39
<< labels >>
rlabel m2contact 2 64 2 64 1 enb
rlabel m2contact 18 45 18 45 1 d
rlabel m2contact 10 37 10 37 1 en
rlabel metal1 -1 0 -1 0 2 Gnd!
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel m2contact 74 55 74 55 1 phi2b
rlabel m2contact 66 45 66 45 1 phi2
rlabel m2contact 90 35 90 35 1 phi1
rlabel m2contact 106 55 106 55 1 phi1b
rlabel m2contact 130 44 130 44 1 q
<< end >>
