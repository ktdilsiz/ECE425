magic
tech scmos
timestamp 1493149052
<< error_s >>
rect -140 -83 -136 -82
<< metal1 >>
rect -350 151 -12 155
rect -8 151 253 155
rect 257 151 258 155
rect -350 144 -60 148
rect -56 144 221 148
rect 225 144 258 148
rect -350 137 -108 141
rect -104 137 189 141
rect 193 137 258 141
rect -350 130 -156 134
rect -152 130 157 134
rect 161 130 258 134
rect -350 123 -204 127
rect -200 123 125 127
rect 129 123 258 127
rect -350 116 -252 120
rect -248 116 93 120
rect 97 116 258 120
rect -350 109 -300 113
rect -296 109 61 113
rect 65 109 258 113
rect -350 102 -348 106
rect -344 102 -261 106
rect -257 102 20 106
rect 24 102 258 106
<< m2contact >>
rect -12 151 -8 155
rect 253 151 257 155
rect -60 144 -56 148
rect 221 144 225 148
rect -108 137 -104 141
rect 189 137 193 141
rect -156 130 -152 134
rect 157 130 161 134
rect -204 123 -200 127
rect 125 123 129 127
rect -252 116 -248 120
rect 93 116 97 120
rect -300 109 -296 113
rect 61 109 65 113
rect -348 102 -344 106
rect -261 102 -257 106
rect 20 102 24 106
rect -324 -20 -320 -16
rect -316 -89 -312 -85
rect -308 -89 -304 -85
rect -330 -97 -326 -93
rect -243 -203 -239 -199
rect -249 -331 -245 -327
rect -249 -340 -245 -336
<< metal2 >>
rect -355 106 -351 107
rect -355 -62 -351 102
rect -348 49 -344 102
rect -324 -16 -320 62
rect -316 -7 -312 51
rect -300 49 -296 109
rect -261 97 -257 102
rect -308 2 -304 45
rect -316 -85 -312 -20
rect -308 -85 -304 -29
rect -300 -89 -296 -11
rect -289 -25 -285 -2
rect -276 -16 -272 62
rect -268 -7 -264 51
rect -252 49 -248 116
rect -268 -81 -264 -29
rect -260 -35 -256 45
rect -228 -16 -224 62
rect -220 -7 -216 51
rect -204 49 -200 123
rect -308 -215 -304 -89
rect -244 -132 -240 -72
rect -236 -83 -232 -29
rect -211 -34 -207 45
rect -197 -25 -193 41
rect -180 -16 -176 62
rect -172 -7 -168 51
rect -156 49 -152 130
rect -160 41 -159 45
rect -211 -39 -207 -38
rect -220 -81 -216 -39
rect -188 -83 -184 -29
rect -163 -34 -159 41
rect -149 -25 -145 41
rect -132 -16 -128 62
rect -124 -7 -120 51
rect -108 49 -104 137
rect -112 41 -111 45
rect -172 -81 -168 -38
rect -163 -39 -159 -38
rect -140 -83 -136 -29
rect -115 -34 -111 41
rect -101 -25 -97 41
rect -84 -16 -80 62
rect -76 -7 -72 51
rect -60 49 -56 144
rect -64 41 -63 45
rect -124 -81 -120 -38
rect -115 -39 -111 -38
rect -92 -83 -88 -29
rect -67 -34 -63 41
rect -53 -25 -49 41
rect -36 -16 -32 62
rect -28 -7 -24 51
rect -12 49 -8 151
rect 12 -16 16 62
rect 20 47 24 102
rect 61 64 65 109
rect 93 64 97 116
rect 125 64 129 123
rect 157 64 161 130
rect 189 64 193 137
rect 221 64 225 144
rect 253 64 257 151
rect -53 -30 -49 -29
rect -76 -81 -72 -38
rect -67 -39 -63 -38
rect -44 -83 -40 -29
rect -28 -81 -24 -38
rect 4 -83 8 -38
rect 20 -81 24 39
rect 28 -51 32 45
rect 36 -25 40 45
rect 52 -16 56 37
rect 36 -30 40 -29
rect 52 -39 56 -33
rect 68 -34 72 45
rect 84 -16 88 37
rect 28 -56 32 -55
rect 52 -43 56 -42
rect 52 -83 56 -47
rect 100 -43 104 45
rect 116 -16 120 37
rect 100 -48 104 -47
rect 68 -81 72 -56
rect 100 -83 104 -56
rect 116 -81 120 -29
rect 132 -51 136 45
rect 148 -16 152 37
rect 164 -25 168 45
rect 180 -16 184 37
rect 148 -83 152 -29
rect 164 -81 168 -46
rect 196 -83 200 45
rect 212 -16 216 37
rect 228 -25 232 45
rect 244 -16 248 37
rect 212 -81 216 -56
rect 244 -83 248 -29
rect -228 -117 -224 -85
rect -180 -131 -176 -85
rect -204 -132 -200 -131
rect -204 -195 -200 -136
rect -172 -211 -168 -121
rect -308 -354 -304 -219
rect -212 -325 -208 -316
rect -148 -321 -144 -202
rect -140 -213 -136 -90
rect -84 -86 -80 -85
rect -36 -86 -32 -85
rect 12 -86 16 -85
rect 60 -86 64 -85
rect 108 -86 112 -85
rect 156 -86 160 -85
rect 204 -86 208 -85
rect 252 -86 256 -85
rect -132 -117 -128 -89
rect -124 -211 -120 -135
rect -92 -213 -88 -90
rect -84 -131 -80 -90
rect -76 -211 -72 -121
rect -44 -213 -40 -90
rect -36 -117 -32 -90
rect -28 -211 -24 -135
rect 4 -213 8 -90
rect 12 -131 16 -90
rect 20 -211 24 -121
rect 52 -213 56 -90
rect 60 -117 64 -90
rect 68 -211 72 -135
rect 100 -213 104 -90
rect 108 -131 112 -90
rect 116 -211 120 -121
rect 148 -213 152 -90
rect 156 -117 160 -90
rect 164 -131 168 -90
rect 164 -211 168 -135
rect 196 -213 200 -90
rect 204 -131 208 -90
rect 212 -211 216 -121
rect 244 -213 248 -90
rect -84 -216 -80 -215
rect 252 -216 256 -215
rect -196 -333 -192 -331
rect -140 -336 -136 -329
rect -124 -341 -120 -220
rect -100 -328 -96 -316
rect -92 -343 -88 -220
rect -76 -341 -72 -220
rect -44 -343 -40 -220
rect -28 -341 -24 -220
rect 4 -343 8 -220
rect 20 -341 24 -220
rect 52 -343 56 -220
rect 68 -341 72 -220
rect 100 -343 104 -220
rect 116 -341 120 -220
rect 148 -343 152 -220
rect 164 -341 168 -220
rect 196 -343 200 -220
rect 212 -341 216 -220
rect 244 -343 248 -220
rect -172 -354 -168 -345
rect -308 -359 -304 -358
rect -84 -396 -80 -345
rect -36 -396 -32 -345
rect 12 -396 16 -345
rect 60 -396 64 -345
rect 108 -396 112 -345
rect 156 -396 160 -345
rect 204 -396 208 -345
rect 252 -396 256 -345
<< m3contact >>
rect -355 102 -351 106
rect -261 102 -257 106
rect -308 -2 -303 2
rect -289 -2 -285 2
rect -316 -11 -312 -7
rect -300 -11 -296 -7
rect -324 -20 -320 -16
rect -316 -20 -312 -16
rect -355 -66 -351 -62
rect -308 -29 -304 -25
rect -268 -11 -264 -7
rect -276 -20 -272 -16
rect -289 -29 -285 -25
rect -268 -29 -264 -25
rect -275 -66 -271 -62
rect -220 -11 -216 -7
rect -228 -20 -224 -16
rect -260 -39 -256 -35
rect -236 -29 -232 -25
rect -244 -72 -240 -68
rect -330 -97 -326 -93
rect -284 -97 -280 -93
rect -197 41 -193 45
rect -164 41 -160 45
rect -172 -11 -168 -7
rect -180 -20 -176 -16
rect -197 -29 -193 -25
rect -188 -29 -184 -25
rect -220 -39 -216 -35
rect -211 -38 -207 -34
rect -196 -72 -192 -68
rect -149 41 -145 45
rect -116 41 -112 45
rect -124 -11 -120 -7
rect -132 -20 -128 -16
rect -149 -29 -145 -25
rect -140 -29 -136 -25
rect -172 -38 -168 -34
rect -163 -38 -159 -34
rect -148 -72 -144 -68
rect -101 41 -97 45
rect -68 41 -64 45
rect -76 -11 -72 -7
rect -84 -20 -80 -16
rect -101 -29 -97 -25
rect -92 -29 -88 -25
rect -124 -38 -120 -34
rect -115 -38 -111 -34
rect -100 -72 -96 -68
rect -53 41 -49 45
rect -20 41 -16 45
rect -28 -11 -24 -7
rect -36 -20 -32 -16
rect 12 -20 16 -16
rect 20 39 24 44
rect -53 -29 -49 -25
rect -44 -29 -40 -25
rect -76 -38 -72 -34
rect -67 -38 -63 -34
rect -52 -72 -48 -68
rect -28 -38 -24 -34
rect 4 -38 8 -34
rect -4 -72 0 -68
rect 52 -20 56 -16
rect 36 -29 40 -25
rect 84 -20 88 -16
rect 68 -38 72 -34
rect 28 -55 32 -51
rect 52 -47 56 -43
rect 44 -72 48 -68
rect 116 -20 120 -16
rect 100 -47 104 -43
rect 116 -29 120 -25
rect 68 -56 72 -52
rect 100 -56 104 -52
rect 92 -72 96 -68
rect 148 -20 152 -16
rect 180 -20 184 -16
rect 132 -55 136 -51
rect 148 -29 152 -25
rect 164 -29 168 -25
rect 140 -72 144 -68
rect 164 -46 168 -42
rect 188 -72 192 -68
rect 212 -20 216 -16
rect 244 -20 248 -16
rect 228 -29 232 -25
rect 244 -29 248 -25
rect 212 -56 216 -52
rect 236 -72 240 -68
rect -228 -121 -224 -117
rect -140 -90 -136 -85
rect -244 -136 -240 -132
rect -204 -136 -200 -132
rect -180 -135 -176 -131
rect -172 -121 -168 -117
rect -243 -203 -239 -199
rect -188 -203 -184 -199
rect -148 -202 -144 -198
rect -308 -219 -304 -215
rect -220 -219 -216 -215
rect -212 -316 -208 -312
rect -132 -89 -128 -85
rect -132 -121 -128 -117
rect -92 -90 -88 -86
rect -124 -135 -120 -131
rect -100 -202 -96 -198
rect -84 -90 -80 -86
rect -44 -90 -40 -86
rect -84 -135 -80 -131
rect -76 -121 -72 -117
rect -52 -202 -48 -198
rect -36 -90 -32 -86
rect -36 -121 -32 -117
rect 4 -90 8 -86
rect -28 -135 -24 -131
rect -4 -202 0 -198
rect 12 -90 16 -86
rect 52 -90 56 -86
rect 12 -135 16 -131
rect 20 -121 24 -117
rect 44 -202 48 -198
rect 60 -90 64 -86
rect 60 -121 64 -117
rect 100 -90 104 -86
rect 68 -135 72 -131
rect 92 -202 96 -198
rect 108 -90 112 -86
rect 148 -90 152 -86
rect 108 -135 112 -131
rect 116 -121 120 -117
rect 140 -202 144 -198
rect 156 -90 160 -86
rect 156 -121 160 -117
rect 164 -90 168 -86
rect 164 -135 168 -131
rect 196 -90 200 -86
rect 188 -202 192 -198
rect 204 -90 208 -86
rect 244 -90 248 -86
rect 252 -90 256 -86
rect 204 -135 208 -131
rect 212 -121 216 -117
rect 236 -202 240 -198
rect -132 -220 -128 -216
rect -124 -220 -120 -216
rect -156 -325 -152 -321
rect -148 -325 -144 -321
rect -249 -331 -245 -327
rect -196 -331 -192 -327
rect -249 -340 -245 -336
rect -140 -340 -136 -336
rect -92 -220 -88 -216
rect -84 -220 -80 -216
rect -76 -220 -72 -216
rect -100 -316 -96 -312
rect -100 -332 -96 -328
rect -44 -220 -40 -216
rect -36 -220 -32 -216
rect -28 -220 -24 -216
rect -52 -332 -48 -328
rect 4 -220 8 -216
rect 12 -220 16 -216
rect 20 -220 24 -216
rect -4 -332 0 -328
rect 52 -220 56 -216
rect 60 -220 64 -216
rect 68 -220 72 -216
rect 44 -332 48 -328
rect 100 -220 104 -216
rect 108 -220 112 -216
rect 116 -220 120 -216
rect 92 -332 96 -328
rect 148 -220 152 -216
rect 156 -220 160 -216
rect 164 -220 168 -216
rect 140 -332 144 -328
rect 196 -220 200 -216
rect 204 -220 208 -216
rect 212 -220 216 -216
rect 188 -332 192 -328
rect 244 -220 248 -216
rect 252 -220 256 -216
rect 236 -332 240 -328
rect -228 -349 -224 -345
rect -308 -358 -304 -354
rect -172 -358 -168 -354
<< metal3 >>
rect -356 106 -256 107
rect -356 102 -355 106
rect -351 102 -261 106
rect -257 102 -256 106
rect -356 101 -256 102
rect -198 45 -159 46
rect -198 41 -197 45
rect -193 41 -164 45
rect -160 41 -159 45
rect -198 40 -159 41
rect -150 45 -111 46
rect -150 41 -149 45
rect -145 41 -116 45
rect -112 41 -111 45
rect -150 40 -111 41
rect -102 45 -63 46
rect -102 41 -101 45
rect -97 41 -68 45
rect -64 41 -63 45
rect -102 40 -63 41
rect -54 45 -15 46
rect -54 41 -53 45
rect -49 41 -20 45
rect -16 44 25 45
rect -16 41 20 44
rect -54 40 20 41
rect -20 39 20 40
rect 24 39 25 44
rect -20 38 25 39
rect -309 2 -284 3
rect -309 -2 -308 2
rect -303 -2 -289 2
rect -285 -2 -284 2
rect -309 -3 -284 -2
rect -348 -7 17 -6
rect -348 -11 -316 -7
rect -312 -11 -300 -7
rect -296 -11 -268 -7
rect -264 -11 -220 -7
rect -216 -11 -172 -7
rect -168 -11 -124 -7
rect -120 -11 -76 -7
rect -72 -11 -28 -7
rect -24 -11 17 -7
rect -348 -12 17 -11
rect -325 -16 256 -15
rect -325 -20 -324 -16
rect -320 -20 -316 -16
rect -312 -20 -276 -16
rect -272 -20 -228 -16
rect -224 -20 -180 -16
rect -176 -20 -132 -16
rect -128 -20 -84 -16
rect -80 -20 -36 -16
rect -32 -20 12 -16
rect 16 -20 52 -16
rect 56 -20 84 -16
rect 88 -20 116 -16
rect 120 -20 148 -16
rect 152 -20 180 -16
rect 184 -20 212 -16
rect 216 -20 244 -16
rect 248 -20 256 -16
rect -325 -21 256 -20
rect -322 -25 -293 -24
rect -322 -29 -308 -25
rect -304 -29 -293 -25
rect -322 -30 -293 -29
rect -290 -25 -263 -24
rect -290 -29 -289 -25
rect -285 -29 -268 -25
rect -264 -29 -263 -25
rect -290 -30 -263 -29
rect -237 -25 -192 -24
rect -237 -29 -236 -25
rect -232 -29 -197 -25
rect -193 -29 -192 -25
rect -237 -30 -192 -29
rect -189 -25 -144 -24
rect -189 -29 -188 -25
rect -184 -29 -149 -25
rect -145 -29 -144 -25
rect -189 -30 -144 -29
rect -141 -25 -96 -24
rect -141 -29 -140 -25
rect -136 -29 -101 -25
rect -97 -29 -96 -25
rect -141 -30 -96 -29
rect -93 -25 -48 -24
rect -93 -29 -92 -25
rect -88 -29 -53 -25
rect -49 -29 -48 -25
rect -93 -30 -48 -29
rect -45 -25 121 -24
rect -45 -29 -44 -25
rect -40 -29 36 -25
rect 40 -29 116 -25
rect 120 -29 121 -25
rect -45 -30 121 -29
rect 147 -25 169 -24
rect 147 -29 148 -25
rect 152 -29 164 -25
rect 168 -29 169 -25
rect 147 -30 169 -29
rect 227 -25 249 -24
rect 227 -29 228 -25
rect 232 -29 244 -25
rect 248 -29 249 -25
rect 227 -30 249 -29
rect -212 -34 -167 -33
rect -261 -35 -215 -34
rect -261 -39 -260 -35
rect -256 -39 -220 -35
rect -216 -39 -215 -35
rect -212 -38 -211 -34
rect -207 -38 -172 -34
rect -168 -38 -167 -34
rect -212 -39 -167 -38
rect -164 -34 -119 -33
rect -164 -38 -163 -34
rect -159 -38 -124 -34
rect -120 -38 -119 -34
rect -164 -39 -119 -38
rect -116 -34 -71 -33
rect -116 -38 -115 -34
rect -111 -38 -76 -34
rect -72 -38 -71 -34
rect -116 -39 -71 -38
rect -68 -34 -23 -33
rect -68 -38 -67 -34
rect -63 -38 -28 -34
rect -24 -38 -23 -34
rect -68 -39 -23 -38
rect 3 -34 36 -33
rect 3 -38 4 -34
rect 8 -38 36 -34
rect 3 -39 36 -38
rect 40 -34 73 -33
rect 40 -38 68 -34
rect 72 -38 73 -34
rect 40 -39 73 -38
rect -261 -40 -215 -39
rect 105 -42 169 -41
rect 51 -43 164 -42
rect 51 -47 52 -43
rect 56 -47 100 -43
rect 104 -46 164 -43
rect 168 -46 169 -42
rect 104 -47 169 -46
rect 51 -48 105 -47
rect 27 -51 41 -50
rect 131 -51 138 -50
rect 27 -55 28 -51
rect 32 -52 73 -51
rect 32 -55 68 -52
rect 27 -56 68 -55
rect 72 -56 73 -52
rect 67 -57 73 -56
rect 99 -52 132 -51
rect 99 -56 100 -52
rect 104 -55 132 -52
rect 136 -52 217 -51
rect 136 -55 212 -52
rect 104 -56 212 -55
rect 216 -56 217 -52
rect 99 -57 217 -56
rect -356 -62 -262 -61
rect -356 -66 -355 -62
rect -351 -66 -275 -62
rect -271 -66 -262 -62
rect -356 -67 -262 -66
rect -246 -68 241 -67
rect -246 -72 -244 -68
rect -240 -72 -196 -68
rect -192 -72 -148 -68
rect -144 -72 -100 -68
rect -96 -72 -52 -68
rect -48 -72 -4 -68
rect 0 -72 44 -68
rect 48 -72 92 -68
rect 96 -72 140 -68
rect 144 -72 188 -68
rect 192 -72 236 -68
rect 240 -72 241 -68
rect -246 -73 241 -72
rect -141 -85 -127 -84
rect -141 -90 -140 -85
rect -136 -89 -132 -85
rect -128 -89 -127 -85
rect -136 -90 -127 -89
rect -141 -91 -127 -90
rect -93 -86 -79 -85
rect -93 -90 -92 -86
rect -88 -90 -84 -86
rect -80 -90 -79 -86
rect -93 -91 -79 -90
rect -45 -86 -31 -85
rect -45 -90 -44 -86
rect -40 -90 -36 -86
rect -32 -90 -31 -86
rect -45 -91 -31 -90
rect 3 -86 17 -85
rect 3 -90 4 -86
rect 8 -90 12 -86
rect 16 -90 17 -86
rect 3 -91 17 -90
rect 51 -86 65 -85
rect 51 -90 52 -86
rect 56 -90 60 -86
rect 64 -90 65 -86
rect 51 -91 65 -90
rect 99 -86 114 -85
rect 99 -90 100 -86
rect 104 -90 108 -86
rect 112 -90 114 -86
rect 99 -91 114 -90
rect 147 -86 169 -85
rect 147 -90 148 -86
rect 152 -90 156 -86
rect 160 -90 164 -86
rect 168 -90 169 -86
rect 147 -91 169 -90
rect 195 -86 209 -85
rect 195 -90 196 -86
rect 200 -90 204 -86
rect 208 -90 209 -86
rect 195 -91 209 -90
rect 243 -86 257 -85
rect 243 -90 244 -86
rect 248 -90 252 -86
rect 256 -90 257 -86
rect 243 -91 257 -90
rect -331 -93 -279 -92
rect -331 -97 -330 -93
rect -326 -97 -284 -93
rect -280 -97 -279 -93
rect -331 -98 -279 -97
rect -229 -117 -167 -116
rect -229 -121 -228 -117
rect -224 -121 -172 -117
rect -168 -121 -167 -117
rect -229 -122 -167 -121
rect -133 -117 -71 -116
rect -133 -121 -132 -117
rect -128 -121 -76 -117
rect -72 -121 -71 -117
rect -133 -122 -71 -121
rect -37 -117 25 -116
rect -37 -121 -36 -117
rect -32 -121 20 -117
rect 24 -121 25 -117
rect -37 -122 25 -121
rect 59 -117 121 -116
rect 59 -121 60 -117
rect 64 -121 116 -117
rect 120 -121 121 -117
rect 59 -122 121 -121
rect 155 -117 217 -116
rect 155 -121 156 -117
rect 160 -121 212 -117
rect 216 -121 217 -117
rect 155 -122 217 -121
rect -181 -131 -119 -130
rect -245 -132 -199 -131
rect -245 -136 -244 -132
rect -240 -136 -204 -132
rect -200 -136 -199 -132
rect -181 -135 -180 -131
rect -176 -135 -124 -131
rect -120 -135 -119 -131
rect -181 -136 -119 -135
rect -85 -131 -23 -130
rect -85 -135 -84 -131
rect -80 -135 -28 -131
rect -24 -135 -23 -131
rect -85 -136 -23 -135
rect 11 -131 73 -130
rect 11 -135 12 -131
rect 16 -135 68 -131
rect 72 -135 73 -131
rect 11 -136 73 -135
rect 107 -131 169 -130
rect 107 -135 108 -131
rect 112 -135 164 -131
rect 168 -135 169 -131
rect 107 -136 169 -135
rect 203 -131 250 -130
rect 203 -135 204 -131
rect 208 -135 250 -131
rect 203 -136 250 -135
rect -245 -137 -199 -136
rect -149 -198 241 -197
rect -244 -199 -183 -198
rect -244 -203 -243 -199
rect -239 -203 -188 -199
rect -184 -203 -183 -199
rect -149 -202 -148 -198
rect -144 -202 -100 -198
rect -96 -202 -52 -198
rect -48 -202 -4 -198
rect 0 -202 44 -198
rect 48 -202 92 -198
rect 96 -202 140 -198
rect 144 -202 188 -198
rect 192 -202 236 -198
rect 240 -202 241 -198
rect -149 -203 241 -202
rect -244 -204 -183 -203
rect -309 -215 -215 -214
rect -309 -219 -308 -215
rect -304 -219 -220 -215
rect -216 -219 -215 -215
rect -309 -220 -215 -219
rect -133 -216 -119 -215
rect -133 -220 -132 -216
rect -128 -220 -124 -216
rect -120 -220 -119 -216
rect -133 -221 -119 -220
rect -93 -216 -71 -215
rect -93 -220 -92 -216
rect -88 -220 -84 -216
rect -80 -220 -76 -216
rect -72 -220 -71 -216
rect -93 -221 -71 -220
rect -45 -216 -23 -215
rect -45 -220 -44 -216
rect -40 -220 -36 -216
rect -32 -220 -28 -216
rect -24 -220 -23 -216
rect -45 -221 -23 -220
rect 3 -216 25 -215
rect 3 -220 4 -216
rect 8 -220 12 -216
rect 16 -220 20 -216
rect 24 -220 25 -216
rect 3 -221 25 -220
rect 51 -216 73 -215
rect 51 -220 52 -216
rect 56 -220 60 -216
rect 64 -220 68 -216
rect 72 -220 73 -216
rect 51 -221 73 -220
rect 99 -216 121 -215
rect 99 -220 100 -216
rect 104 -220 108 -216
rect 112 -220 116 -216
rect 120 -220 121 -216
rect 99 -221 121 -220
rect 147 -216 169 -215
rect 147 -220 148 -216
rect 152 -220 156 -216
rect 160 -220 164 -216
rect 168 -220 169 -216
rect 147 -221 169 -220
rect 195 -216 217 -215
rect 195 -220 196 -216
rect 200 -220 204 -216
rect 208 -220 212 -216
rect 216 -220 217 -216
rect 195 -221 217 -220
rect 243 -216 257 -215
rect 243 -220 244 -216
rect 248 -220 252 -216
rect 256 -220 257 -216
rect 243 -221 257 -220
rect -213 -312 -95 -311
rect -213 -316 -212 -312
rect -208 -316 -100 -312
rect -96 -316 -95 -312
rect -213 -317 -95 -316
rect -157 -321 -143 -320
rect -157 -325 -156 -321
rect -152 -325 -148 -321
rect -144 -325 -143 -321
rect -157 -326 -143 -325
rect -250 -327 -191 -326
rect -250 -331 -249 -327
rect -245 -331 -196 -327
rect -192 -331 -191 -327
rect -250 -332 -191 -331
rect -101 -328 241 -327
rect -101 -332 -100 -328
rect -96 -332 -52 -328
rect -48 -332 -4 -328
rect 0 -332 44 -328
rect 48 -332 92 -328
rect 96 -332 140 -328
rect 144 -332 188 -328
rect 192 -332 236 -328
rect 240 -332 241 -328
rect -101 -333 241 -332
rect -250 -336 -135 -335
rect -250 -340 -249 -336
rect -245 -340 -140 -336
rect -136 -340 -135 -336
rect -250 -341 -135 -340
rect -249 -345 -223 -344
rect -249 -349 -228 -345
rect -224 -349 -223 -345
rect -249 -350 -223 -349
rect -249 -353 -243 -350
rect -309 -354 -167 -353
rect -309 -358 -308 -354
rect -304 -358 -172 -354
rect -168 -358 -167 -354
rect -309 -359 -167 -358
use mux2_dp_1x  mux2_dp_1x_0
timestamp 1484435125
transform 1 0 -348 0 1 3
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_1
timestamp 1484435125
transform 1 0 -300 0 1 3
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_2
timestamp 1484435125
transform 1 0 -252 0 1 3
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_3
timestamp 1484435125
transform 1 0 -204 0 1 3
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_4
timestamp 1484435125
transform 1 0 -156 0 1 3
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_5
timestamp 1484435125
transform 1 0 -108 0 1 3
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_6
timestamp 1484435125
transform 1 0 -60 0 1 3
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_7
timestamp 1484435125
transform 1 0 -12 0 1 3
box -6 -4 50 96
use and2_1x  and2_1x_0
timestamp 1484419738
transform 1 0 36 0 1 3
box -6 -4 34 96
use and2_1x  and2_1x_1
timestamp 1484419738
transform 1 0 68 0 1 3
box -6 -4 34 96
use and2_1x  and2_1x_2
timestamp 1484419738
transform 1 0 100 0 1 3
box -6 -4 34 96
use and2_1x  and2_1x_3
timestamp 1484419738
transform 1 0 132 0 1 3
box -6 -4 34 96
use and2_1x  and2_1x_4
timestamp 1484419738
transform 1 0 164 0 1 3
box -6 -4 34 96
use and2_1x  and2_1x_5
timestamp 1484419738
transform 1 0 196 0 1 3
box -6 -4 34 96
use and2_1x  and2_1x_6
timestamp 1484419738
transform 1 0 228 0 1 3
box -6 -4 34 96
use inv_1x  inv_1x_0
timestamp 1484418501
transform 1 0 -316 0 1 -127
box -6 -4 18 96
use and2_1x  and2_1x_7
timestamp 1484419738
transform 1 0 -300 0 1 -127
box -6 -4 34 96
use mux2_dp_1x  mux2_dp_1x_20
timestamp 1484435125
transform 1 0 -268 0 1 -127
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_17
timestamp 1484435125
transform 1 0 -220 0 1 -127
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_16
timestamp 1484435125
transform 1 0 -172 0 1 -127
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_15
timestamp 1484435125
transform 1 0 -124 0 1 -127
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_14
timestamp 1484435125
transform 1 0 -76 0 1 -127
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_13
timestamp 1484435125
transform 1 0 -28 0 1 -127
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_12
timestamp 1484435125
transform 1 0 20 0 1 -127
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_11
timestamp 1484435125
transform 1 0 68 0 1 -127
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_10
timestamp 1484435125
transform 1 0 116 0 1 -127
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_9
timestamp 1484435125
transform 1 0 164 0 1 -127
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_8
timestamp 1484435125
transform 1 0 212 0 1 -127
box -6 -4 50 96
use xor2_1x  xor2_1x_0
timestamp 1492273518
transform 1 0 -228 0 1 -257
box -6 -4 58 96
use mux2_dp_1x  mux2_dp_1x_27
timestamp 1484435125
transform 1 0 -172 0 1 -257
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_26
timestamp 1484435125
transform 1 0 -124 0 1 -257
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_25
timestamp 1484435125
transform 1 0 -76 0 1 -257
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_24
timestamp 1484435125
transform 1 0 -28 0 1 -257
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_23
timestamp 1484435125
transform 1 0 20 0 1 -257
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_22
timestamp 1484435125
transform 1 0 68 0 1 -257
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_21
timestamp 1484435125
transform 1 0 116 0 1 -257
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_19
timestamp 1484435125
transform 1 0 164 0 1 -257
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_18
timestamp 1484435125
transform 1 0 212 0 1 -257
box -6 -4 50 96
use xor2_1x  xor2_1x_2
timestamp 1492273518
transform 1 0 -236 0 1 -387
box -6 -4 58 96
use xor2_1x  xor2_1x_1
timestamp 1492273518
transform 1 0 -180 0 1 -387
box -6 -4 58 96
use mux2_dp_1x  mux2_dp_1x_35
timestamp 1484435125
transform 1 0 -124 0 1 -387
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_34
timestamp 1484435125
transform 1 0 -76 0 1 -387
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_33
timestamp 1484435125
transform 1 0 -28 0 1 -387
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_32
timestamp 1484435125
transform 1 0 20 0 1 -387
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_31
timestamp 1484435125
transform 1 0 68 0 1 -387
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_30
timestamp 1484435125
transform 1 0 116 0 1 -387
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_29
timestamp 1484435125
transform 1 0 164 0 1 -387
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_28
timestamp 1484435125
transform 1 0 212 0 1 -387
box -6 -4 50 96
<< labels >>
rlabel metal1 -348 111 -348 111 1 a6
rlabel metal1 -348 118 -348 118 1 a5
rlabel metal1 -348 125 -348 125 1 a4
rlabel metal1 -348 132 -348 132 1 a3
rlabel metal1 -348 139 -348 139 1 a2
rlabel metal1 -348 146 -348 146 1 a1
rlabel metal1 -348 153 -348 153 5 a0
rlabel m3contact -328 -95 -328 -95 1 arith
rlabel metal3 -320 -27 -320 -27 1 rightb
rlabel metal3 -320 -9 -320 -9 1 arithAndRight
rlabel metal1 -348 104 -348 104 1 a7
rlabel metal3 -241 -217 -241 -217 1 rightinverse
rlabel metal3 -247 -356 -247 -356 1 rightinverse
rlabel metal3 -247 -347 -247 -347 1 rightinverse
rlabel m3contact -322 -18 -322 -18 1 right
rlabel metal2 -82 -394 -82 -394 1 Y7
rlabel metal2 -34 -394 -34 -394 1 Y6
rlabel metal2 14 -394 14 -394 1 Y5
rlabel metal2 62 -394 62 -394 1 Y4
rlabel metal2 110 -394 110 -394 1 Y3
rlabel metal2 158 -394 158 -394 1 Y2
rlabel metal2 206 -394 206 -394 1 Y1
rlabel metal2 254 -394 254 -394 1 Y0
rlabel m3contact -241 -201 -241 -201 1 Shamt_2
rlabel m3contact -247 -329 -247 -329 1 Shamt_0
rlabel m3contact -247 -338 -247 -338 1 Shamt_1
rlabel metal2 -306 42 -306 42 1 Z14
rlabel metal2 -258 42 -258 42 1 Z13
rlabel metal2 -210 42 -210 42 1 Z12
rlabel m3contact -162 42 -162 42 1 Z11
rlabel m3contact -114 42 -114 42 1 Z10
rlabel m3contact -66 42 -66 42 1 Z09
rlabel m3contact -18 42 -18 42 1 Z08
rlabel metal2 30 42 30 42 1 Z07
rlabel metal2 38 42 38 42 1 Z06
rlabel metal2 70 42 70 42 1 Z05
rlabel metal2 102 42 102 42 1 Z04
rlabel metal2 134 42 134 42 1 Z03
rlabel metal2 166 42 166 42 1 Z02
rlabel metal2 198 42 198 42 1 Z01
rlabel metal2 230 42 230 42 1 Z00
<< end >>
