magic
tech scmos
timestamp 1486497882
use and2_1x  and2_1x_0
array 0 0 40 0 7 110
timestamp 1484419738
transform 1 0 6 0 1 4
box -6 -4 34 96
<< end >>
