magic
tech scmos
timestamp 1494281060
<< metal1 >>
rect 3961 3850 4007 3851
rect 3965 3846 4007 3850
rect 3961 3845 4007 3846
rect 3968 3550 4006 3551
rect 3972 3546 4006 3550
rect 3968 3544 4006 3546
rect 2904 3275 2960 3276
rect 2904 3271 3965 3275
rect 2904 3267 3961 3271
rect 2904 3262 3965 3267
rect 2904 3261 2960 3262
rect 2904 3212 2916 3261
rect 1105 3200 1208 3207
rect 1105 3176 1109 3200
rect 1067 3086 1074 3094
rect 1067 2991 1071 3086
rect 1119 3080 1124 3200
rect 2205 3198 2916 3212
rect 2920 3237 2935 3239
rect 2920 3235 2941 3237
rect 2920 3230 2935 3235
rect 2940 3230 2941 3235
rect 2920 3228 2941 3230
rect 2920 3185 2935 3228
rect 2176 3173 2935 3185
rect 1104 3074 1124 3080
rect 2920 3030 2935 3173
rect 2929 3021 2935 3030
rect 2945 2998 2960 3261
rect 2964 3235 3972 3237
rect 2964 3230 2965 3235
rect 2970 3231 3968 3235
rect 2970 3230 3972 3231
rect 2964 3228 3972 3230
rect 3815 3134 3965 3135
rect 3815 3130 3961 3134
rect 3815 3127 3965 3130
rect 3815 3043 3972 3045
rect 3815 3039 3968 3043
rect 3815 3037 3972 3039
rect 3815 3003 3965 3005
rect 3815 2999 3961 3003
rect 3815 2997 3965 2999
rect 1067 2990 1074 2991
rect 1067 2989 1076 2990
rect 1067 2985 1069 2989
rect 1073 2985 1076 2989
rect 1067 2984 1076 2985
rect 1067 2983 1074 2984
rect 3815 2913 3972 2915
rect 3815 2909 3968 2913
rect 3815 2907 3972 2909
rect 3815 2873 3965 2875
rect 3815 2869 3961 2873
rect 3815 2867 3965 2869
rect 3815 2783 3972 2785
rect 3815 2779 3968 2783
rect 3815 2777 3972 2779
rect 3815 2743 3965 2745
rect 3815 2739 3961 2743
rect 3815 2737 3965 2739
rect 3815 2654 3972 2655
rect 3815 2650 3968 2654
rect 3815 2647 3972 2650
rect 3910 2484 3965 2486
rect 3910 2480 3961 2484
rect 3910 2478 3965 2480
rect 3958 2394 3972 2396
rect 3958 2390 3968 2394
rect 3958 2388 3972 2390
rect 3910 2375 3965 2376
rect 3910 2371 3961 2375
rect 3910 2368 3965 2371
rect 3958 2284 3972 2286
rect 3958 2280 3968 2284
rect 3958 2278 3972 2280
rect 3910 2264 3965 2266
rect 3910 2260 3961 2264
rect 3910 2258 3965 2260
rect 3958 2174 3972 2176
rect 3958 2170 3968 2174
rect 3958 2168 3972 2170
rect 3910 2155 3965 2156
rect 3910 2151 3961 2155
rect 3910 2148 3965 2151
rect 3958 2064 3972 2066
rect 3958 2060 3968 2064
rect 3958 2058 3972 2060
rect 3910 2044 3965 2046
rect 3910 2040 3961 2044
rect 3910 2038 3965 2040
rect 3958 1954 3972 1956
rect 3958 1950 3968 1954
rect 3958 1948 3972 1950
rect 3910 1934 3965 1936
rect 3910 1930 3961 1934
rect 3910 1928 3965 1930
rect 3958 1844 3972 1846
rect 3958 1840 3968 1844
rect 3958 1838 3972 1840
rect 3910 1824 3965 1826
rect 3910 1820 3961 1824
rect 3910 1818 3965 1820
rect 3958 1734 3972 1736
rect 3958 1730 3968 1734
rect 3958 1728 3972 1730
rect 3910 1715 3965 1716
rect 3910 1711 3961 1715
rect 3910 1708 3965 1711
rect 3958 1624 3972 1626
rect 3958 1620 3968 1624
rect 3958 1618 3972 1620
rect 3910 1604 3965 1606
rect 3910 1600 3961 1604
rect 3910 1598 3965 1600
rect 3958 1514 3972 1516
rect 3958 1510 3968 1514
rect 3958 1508 3972 1510
rect 3910 1494 3965 1496
rect 3910 1490 3961 1494
rect 3910 1488 3965 1490
rect 3958 1404 3972 1406
rect 3958 1400 3968 1404
rect 3958 1398 3972 1400
rect 3910 1384 3965 1386
rect 3910 1380 3961 1384
rect 3910 1378 3965 1380
rect 3958 1294 3972 1296
rect 3958 1290 3968 1294
rect 3958 1288 3972 1290
rect 3910 1274 3965 1276
rect 3910 1270 3961 1274
rect 3910 1268 3965 1270
rect 3958 1184 3972 1186
rect 3958 1180 3968 1184
rect 3958 1178 3972 1180
<< m2contact >>
rect 3961 3846 3965 3850
rect 3968 3546 3972 3550
rect 3961 3267 3965 3271
rect 2935 3230 2940 3235
rect 2920 3021 2929 3030
rect 2965 3230 2970 3235
rect 3968 3231 3972 3235
rect 3961 3130 3965 3134
rect 3968 3039 3972 3043
rect 3961 2999 3965 3003
rect 1069 2985 1073 2989
rect 3968 2909 3972 2913
rect 3961 2869 3965 2873
rect 3968 2779 3972 2783
rect 3961 2739 3965 2743
rect 3968 2650 3972 2654
rect 3961 2480 3965 2484
rect 3968 2390 3972 2394
rect 3961 2371 3965 2375
rect 3968 2280 3972 2284
rect 3961 2260 3965 2264
rect 3968 2170 3972 2174
rect 3961 2151 3965 2155
rect 3968 2060 3972 2064
rect 3961 2040 3965 2044
rect 3968 1950 3972 1954
rect 3961 1930 3965 1934
rect 3968 1840 3972 1844
rect 3961 1820 3965 1824
rect 3968 1730 3972 1734
rect 3961 1711 3965 1715
rect 3968 1620 3972 1624
rect 3961 1600 3965 1604
rect 3968 1510 3972 1514
rect 3961 1490 3965 1494
rect 3968 1400 3972 1404
rect 3961 1380 3965 1384
rect 3968 1290 3972 1294
rect 3961 1270 3965 1274
rect 3968 1180 3972 1184
<< metal2 >>
rect 1259 3998 1263 4000
rect 992 3359 1013 3363
rect 1008 3070 1012 3359
rect 1016 3077 1020 3992
rect 3961 3850 3965 3962
rect 3961 3271 3965 3846
rect 2933 3235 2990 3238
rect 2933 3230 2935 3235
rect 2940 3230 2965 3235
rect 2970 3230 2990 3235
rect 2933 3228 2990 3230
rect 3961 3134 3965 3267
rect 1016 3073 1028 3077
rect 1008 3066 1021 3070
rect 992 3059 1014 3063
rect 1010 2770 1014 3059
rect 1017 2777 1021 3066
rect 1024 2784 1028 3073
rect 2920 3030 2935 3032
rect 2929 3021 2935 3030
rect 2920 2992 2935 3021
rect 3961 3003 3965 3130
rect 3961 2873 3965 2999
rect 1024 2780 1032 2784
rect 1017 2773 1025 2777
rect 1010 2766 1018 2770
rect 993 2759 1011 2763
rect 1007 2471 1011 2759
rect 1014 2478 1018 2766
rect 1021 2485 1025 2773
rect 1028 2498 1032 2780
rect 3961 2743 3965 2869
rect 1035 2498 1039 2502
rect 1028 2494 1039 2498
rect 1021 2481 1032 2485
rect 1014 2474 1025 2478
rect 1007 2467 1018 2471
rect 992 2459 1006 2463
rect 1014 2456 1018 2467
rect 1006 2452 1018 2456
rect 1006 2170 1010 2452
rect 1006 2166 1016 2170
rect 992 2159 1005 2163
rect 1012 2156 1016 2166
rect 1006 2152 1016 2156
rect 1006 1871 1010 2152
rect 1021 1925 1025 2474
rect 1028 2035 1032 2481
rect 1035 2476 1039 2494
rect 1195 2490 1199 2556
rect 3961 2484 3965 2739
rect 1175 2459 1176 2463
rect 1172 2388 1176 2459
rect 1171 2376 1175 2388
rect 1028 2030 1030 2035
rect 1028 2027 1032 2030
rect 1028 2023 1034 2027
rect 1021 1920 1022 1925
rect 1021 1879 1025 1920
rect 1021 1875 1027 1879
rect 1006 1867 1019 1871
rect 993 1859 1007 1863
rect 1015 1815 1019 1867
rect 1015 1807 1019 1810
rect 1172 1705 1176 2376
rect 3961 2375 3965 2480
rect 3961 2264 3965 2371
rect 1172 1699 1176 1700
rect 1195 1595 1199 2159
rect 3961 2155 3965 2260
rect 3961 2044 3965 2151
rect 3961 1934 3965 2040
rect 1203 1485 1207 1859
rect 3961 1824 3965 1930
rect 3961 1715 3965 1820
rect 3961 1604 3965 1711
rect 3961 1494 3965 1600
rect 3961 1384 3965 1490
rect 992 1346 1005 1350
rect 3961 1274 3965 1380
rect 1203 1051 1207 1259
rect 3961 1150 3965 1270
rect 3968 3550 3975 3551
rect 3972 3546 3975 3550
rect 3968 3544 3975 3546
rect 3968 3235 3972 3544
rect 3968 3043 3972 3231
rect 3968 2913 3972 3039
rect 3968 2783 3972 2909
rect 3968 2654 3972 2779
rect 3968 2394 3972 2650
rect 3968 2284 3972 2390
rect 3968 2174 3972 2280
rect 3968 2064 3972 2170
rect 3968 1954 3972 2060
rect 3968 1844 3972 1950
rect 3968 1734 3972 1840
rect 3968 1624 3972 1730
rect 3968 1514 3972 1620
rect 3968 1404 3972 1510
rect 3968 1294 3972 1400
rect 3968 1184 3972 1290
rect 3968 1150 3972 1180
rect 992 1046 1011 1050
<< m3contact >>
rect 1257 4000 1266 4009
rect 1016 3992 1021 3997
rect 991 3957 1000 3966
rect 991 3657 1000 3666
rect 1069 2985 1073 2989
rect 1231 2985 1236 2990
rect 1006 2459 1011 2464
rect 1005 2159 1009 2163
rect 1187 2487 1191 2491
rect 1035 2471 1040 2476
rect 1170 2459 1175 2464
rect 1030 2030 1035 2035
rect 1022 1920 1027 1925
rect 1007 1859 1012 1864
rect 1015 1810 1020 1815
rect 1195 2159 1200 2164
rect 1172 1700 1177 1705
rect 1203 1859 1208 1864
rect 1195 1590 1200 1595
rect 1203 1480 1208 1485
rect 1005 1346 1010 1351
rect 1203 1259 1208 1264
rect 1203 1046 1208 1051
<< metal3 >>
rect 1256 4009 1267 4010
rect 1256 4007 1257 4009
rect 1046 4001 1257 4007
rect 1015 3997 1022 3998
rect 1046 3997 1052 4001
rect 1256 4000 1257 4001
rect 1266 4000 1267 4009
rect 1256 3999 1267 4000
rect 1015 3992 1016 3997
rect 1021 3992 1052 3997
rect 1015 3991 1052 3992
rect 990 3966 1001 3967
rect 990 3957 991 3966
rect 1000 3964 1001 3966
rect 1000 3958 1021 3964
rect 1000 3957 1001 3958
rect 990 3956 1001 3957
rect 990 3666 1001 3667
rect 990 3657 991 3666
rect 1000 3664 1001 3666
rect 1000 3658 1012 3664
rect 1000 3657 1001 3658
rect 990 3656 1001 3657
rect 1006 2492 1012 3658
rect 1015 2557 1021 3958
rect 1230 2990 1237 2991
rect 1068 2989 1231 2990
rect 1068 2985 1069 2989
rect 1073 2985 1231 2989
rect 1236 2985 1237 2990
rect 1068 2984 1237 2985
rect 1015 2551 1200 2557
rect 1006 2491 1192 2492
rect 1006 2487 1187 2491
rect 1191 2487 1192 2491
rect 1006 2486 1192 2487
rect 1034 2476 1041 2477
rect 1034 2471 1035 2476
rect 1040 2471 1184 2476
rect 1034 2470 1184 2471
rect 1005 2464 1012 2465
rect 1169 2464 1176 2465
rect 1005 2459 1006 2464
rect 1011 2459 1170 2464
rect 1175 2459 1178 2464
rect 1005 2458 1178 2459
rect 1178 2379 1179 2380
rect 1194 2164 1201 2165
rect 1004 2163 1195 2164
rect 1004 2159 1005 2163
rect 1009 2159 1195 2163
rect 1200 2159 1212 2164
rect 1004 2158 1212 2159
rect 1029 2035 1036 2036
rect 1027 2030 1030 2035
rect 1035 2030 1202 2035
rect 1027 2029 1202 2030
rect 1021 1925 1028 1926
rect 1021 1920 1022 1925
rect 1027 1920 1202 1925
rect 1021 1919 1202 1920
rect 1006 1864 1013 1865
rect 1202 1864 1209 1865
rect 1006 1859 1007 1864
rect 1012 1859 1203 1864
rect 1208 1859 1212 1864
rect 1006 1858 1212 1859
rect 1014 1815 1021 1816
rect 1014 1810 1015 1815
rect 1020 1810 1202 1815
rect 1014 1809 1202 1810
rect 1171 1705 1178 1706
rect 1171 1700 1172 1705
rect 1177 1700 1202 1705
rect 1171 1699 1202 1700
rect 1194 1595 1201 1596
rect 1194 1590 1195 1595
rect 1200 1590 1202 1595
rect 1194 1589 1202 1590
rect 1202 1485 1209 1486
rect 1202 1480 1203 1485
rect 1208 1480 1209 1485
rect 1202 1479 1209 1480
rect 1132 1359 1203 1365
rect 1004 1351 1011 1352
rect 1132 1351 1138 1359
rect 1004 1346 1005 1351
rect 1010 1346 1138 1351
rect 1004 1345 1138 1346
rect 1202 1264 1209 1265
rect 1202 1259 1203 1264
rect 1208 1259 1209 1264
rect 1202 1258 1209 1259
rect 1194 1249 1205 1255
rect 1187 1239 1206 1245
rect 1202 1051 1209 1052
rect 1005 1046 1203 1051
rect 1208 1046 1211 1051
rect 1005 1045 1211 1046
<< m2p >>
rect 1002 1859 1003 1863
use PADFC  PADFC_0
timestamp 949001400
transform 1 0 0 0 1 4000
box 327 -3 1003 673
use PADINC  reset
timestamp 1084294328
transform 1 0 1000 0 1 4000
box -6 -3 303 1000
use PADOUT  adr0
timestamp 1084294529
transform 1 0 1300 0 1 4000
box -6 -3 303 1000
use PADOUT  adr1
timestamp 1084294529
transform 1 0 1600 0 1 4000
box -6 -3 303 1000
use PADOUT  adr2
timestamp 1084294529
transform 1 0 1900 0 1 4000
box -6 -3 303 1000
use PADOUT  adr3
timestamp 1084294529
transform 1 0 2200 0 1 4000
box -6 -3 303 1000
use PADOUT  adr4
timestamp 1084294529
transform 1 0 2500 0 1 4000
box -6 -3 303 1000
use PADOUT  adr5
timestamp 1084294529
transform 1 0 2800 0 1 4000
box -6 -3 303 1000
use PADOUT  adr6
timestamp 1084294529
transform 1 0 3100 0 1 4000
box -6 -3 303 1000
use PADOUT  adr7
timestamp 1084294529
transform 1 0 3400 0 1 4000
box -6 -3 303 1000
use PADOUT  MemWrite
timestamp 1084294529
transform 1 0 3700 0 1 4000
box -6 -3 303 1000
use PADFC  PADFC_3
timestamp 949001400
transform 0 1 4000 -1 0 5000
box 327 -3 1003 673
use PADINC  ph1
timestamp 1084294328
transform 0 -1 1000 1 0 3700
box -6 -3 303 1000
use PADINC  ph2
timestamp 1084294328
transform 0 -1 1000 1 0 3400
box -6 -3 303 1000
use PADVDD  PADVDD_0
timestamp 1084294447
transform 0 1 4000 -1 0 3997
box -3 -3 303 1000
use PADGND  PADGND_0
timestamp 1084294269
transform 0 1 4000 -1 0 3698
box -3 -3 303 1000
use PADINC  memdata7
timestamp 1084294328
transform 0 -1 1000 1 0 3100
box -6 -3 303 1000
use PADINC  memdata6
timestamp 1084294328
transform 0 -1 1000 1 0 2800
box -6 -3 303 1000
use PADINC  memdata5
timestamp 1084294328
transform 0 -1 1000 1 0 2500
box -6 -3 303 1000
use PADINC  memdata4
timestamp 1084294328
transform 0 -1 1000 1 0 2200
box -6 -3 303 1000
use PADINC  memdata3
timestamp 1084294328
transform 0 -1 1000 1 0 1900
box -6 -3 303 1000
use PADINC  memdata2
timestamp 1084294328
transform 0 -1 1000 1 0 1600
box -6 -3 303 1000
use PADOUT  memdata1
timestamp 1084294529
transform 0 -1 1000 1 0 1300
box -6 -3 303 1000
use datapath  datapath_0
timestamp 1494278851
transform 1 0 1219 0 1 1182
box -168 -32 2739 2085
use PADNC  PADNC_9
timestamp 1084294400
transform 0 1 4000 1 0 3100
box -3 -3 303 1000
use PADNC  PADNC_8
timestamp 1084294400
transform 0 1 4000 1 0 2800
box -3 -3 303 1000
use PADNC  PADNC_7
timestamp 1084294400
transform 0 1 4000 1 0 2500
box -3 -3 303 1000
use PADNC  PADNC_6
timestamp 1084294400
transform 0 1 4000 1 0 2200
box -3 -3 303 1000
use PADNC  PADNC_5
timestamp 1084294400
transform 0 1 4000 1 0 1900
box -3 -3 303 1000
use PADNC  PADNC_4
timestamp 1084294400
transform 0 1 4000 1 0 1600
box -3 -3 303 1000
use PADNC  PADNC_3
timestamp 1084294400
transform 0 1 4000 1 0 1300
box -3 -3 303 1000
use PADOUT  memdata0
timestamp 1084294529
transform 0 -1 1000 1 0 1000
box -6 -3 303 1000
use PADFC  PADFC_2
timestamp 949001400
transform 0 -1 1000 1 0 0
box 327 -3 1003 673
use PADOUT  writedata0
timestamp 1084294529
transform -1 0 1300 0 -1 1000
box -6 -3 303 1000
use PADOUT  writedata1
timestamp 1084294529
transform -1 0 1600 0 -1 1000
box -6 -3 303 1000
use PADOUT  writedata2
timestamp 1084294529
transform -1 0 1900 0 -1 1000
box -6 -3 303 1000
use PADOUT  writedata3
timestamp 1084294529
transform -1 0 2200 0 -1 1000
box -6 -3 303 1000
use PADOUT  writedata4
timestamp 1084294529
transform -1 0 2500 0 -1 1000
box -6 -3 303 1000
use PADOUT  writedata5
timestamp 1084294529
transform -1 0 2800 0 -1 1000
box -6 -3 303 1000
use PADOUT  writedata6
timestamp 1084294529
transform -1 0 3100 0 -1 1000
box -6 -3 303 1000
use PADOUT  writedata7
timestamp 1084294529
transform -1 0 3400 0 -1 1000
box -6 -3 303 1000
use PADNC  PADNC_0
timestamp 1084294400
transform 1 0 3400 0 -1 1000
box -3 -3 303 1000
use PADNC  PADNC_1
timestamp 1084294400
transform 0 1 4000 1 0 1000
box -3 -3 303 1000
use PADFC  PADFC_1
timestamp 949001400
transform -1 0 4998 0 -1 1000
box 327 -3 1003 673
use PADNC  PADNC_2
timestamp 1084294400
transform 1 0 3700 0 -1 1000
box -3 -3 303 1000
<< end >>
