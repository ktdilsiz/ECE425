magic
tech scmos
timestamp 1491245670
<< nwell >>
rect 209 297 497 332
rect -6 53 29 285
rect 29 -8 497 26
<< ntransistor >>
rect 48 179 50 183
rect 56 179 58 183
rect 48 171 50 175
rect 56 171 58 175
rect 40 155 42 159
rect 40 147 42 151
rect 40 131 42 135
rect 56 155 58 159
rect 56 147 58 151
rect 56 131 58 135
rect 48 123 50 127
rect 56 123 58 127
rect 48 107 50 111
rect 56 107 58 111
rect 40 38 42 43
rect 56 38 58 43
rect 80 179 82 183
rect 88 179 90 183
rect 72 171 74 175
rect 72 155 74 159
rect 72 147 74 151
rect 72 131 74 135
rect 88 171 90 175
rect 88 155 90 159
rect 104 179 106 183
rect 104 171 106 175
rect 120 179 122 183
rect 120 171 122 175
rect 112 155 114 159
rect 120 155 122 159
rect 96 147 98 151
rect 104 147 106 151
rect 88 131 90 135
rect 80 123 82 127
rect 88 123 90 127
rect 72 107 74 111
rect 72 38 74 43
rect 88 107 90 111
rect 88 38 90 43
rect 104 131 106 135
rect 104 123 106 127
rect 104 107 106 111
rect 104 38 106 43
rect 120 147 122 151
rect 120 131 122 135
rect 120 123 122 127
rect 120 107 122 111
rect 120 38 122 43
rect 144 275 146 279
rect 144 267 146 271
rect 160 275 162 279
rect 168 275 170 279
rect 160 267 162 271
rect 168 267 170 271
rect 144 251 146 255
rect 152 251 154 255
rect 144 243 146 247
rect 152 243 154 247
rect 144 227 146 231
rect 152 227 154 231
rect 144 219 146 223
rect 152 219 154 223
rect 136 203 138 207
rect 136 195 138 199
rect 136 179 138 183
rect 136 171 138 175
rect 136 155 138 159
rect 136 147 138 151
rect 136 131 138 135
rect 136 123 138 127
rect 136 107 138 111
rect 136 99 138 103
rect 136 83 138 87
rect 136 75 138 79
rect 136 59 138 63
rect 136 38 138 43
rect 192 275 194 279
rect 375 276 379 278
rect 184 267 186 271
rect 176 251 178 255
rect 255 268 259 270
rect 335 268 339 270
rect 192 251 194 255
rect 231 252 235 254
rect 239 252 243 254
rect 351 252 355 254
rect 407 252 411 254
rect 176 243 178 247
rect 184 243 186 247
rect 168 227 170 231
rect 168 219 170 223
rect 160 203 162 207
rect 160 195 162 199
rect 359 244 363 246
rect 375 244 379 246
rect 192 227 194 231
rect 215 228 219 230
rect 407 228 411 230
rect 447 228 451 230
rect 471 228 475 230
rect 184 219 186 223
rect 176 203 178 207
rect 383 220 387 222
rect 423 220 427 222
rect 192 203 194 207
rect 375 204 379 206
rect 399 204 403 206
rect 176 195 178 199
rect 184 195 186 199
rect 160 179 162 183
rect 168 179 170 183
rect 160 171 162 175
rect 168 171 170 175
rect 160 155 162 159
rect 168 155 170 159
rect 160 147 162 151
rect 168 147 170 151
rect 160 131 162 135
rect 168 131 170 135
rect 160 123 162 127
rect 168 123 170 127
rect 160 107 162 111
rect 168 107 170 111
rect 152 99 154 103
rect 152 83 154 87
rect 152 75 154 79
rect 152 59 154 63
rect 152 38 154 43
rect 383 196 387 198
rect 431 196 435 198
rect 455 196 459 198
rect 471 196 475 198
rect 479 196 483 198
rect 192 179 194 183
rect 311 180 315 182
rect 407 180 411 182
rect 447 180 451 182
rect 192 171 194 175
rect 311 172 315 174
rect 407 172 411 174
rect 455 172 459 174
rect 471 172 475 174
rect 184 155 186 159
rect 184 147 186 151
rect 184 131 186 135
rect 184 123 186 127
rect 184 107 186 111
rect 176 99 178 103
rect 311 156 315 158
rect 327 156 331 158
rect 447 156 451 158
rect 455 156 459 158
rect 311 148 315 150
rect 327 148 331 150
rect 447 148 451 150
rect 471 148 475 150
rect 479 148 483 150
rect 311 132 315 134
rect 327 132 331 134
rect 447 132 451 134
rect 479 132 483 134
rect 311 124 315 126
rect 327 124 331 126
rect 455 124 459 126
rect 479 124 483 126
rect 311 108 315 110
rect 327 108 331 110
rect 455 108 459 110
rect 479 108 483 110
rect 192 99 194 103
rect 255 100 259 102
rect 263 100 267 102
rect 327 100 331 102
rect 431 100 435 102
rect 455 100 459 102
rect 176 83 178 87
rect 184 83 186 87
rect 168 75 170 79
rect 168 59 170 63
rect 168 38 170 43
rect 255 84 259 86
rect 279 84 283 86
rect 327 84 331 86
rect 431 84 435 86
rect 471 84 475 86
rect 479 84 483 86
rect 192 75 194 79
rect 255 76 259 78
rect 287 76 291 78
rect 327 76 331 78
rect 431 76 435 78
rect 471 76 475 78
rect 184 59 186 63
rect 184 38 186 43
rect 255 60 259 62
rect 303 60 307 62
rect 327 60 331 62
rect 431 60 435 62
rect 479 60 483 62
rect 220 38 222 43
rect 228 38 230 43
rect 244 38 246 43
rect 252 38 254 43
rect 268 38 270 43
rect 276 38 278 43
rect 292 38 294 43
rect 300 38 302 43
rect 316 38 318 43
rect 324 38 326 43
rect 340 38 342 43
rect 348 38 350 43
rect 364 38 366 43
rect 372 38 374 43
rect 388 38 390 43
rect 396 38 398 43
rect 412 38 414 43
rect 420 38 422 43
rect 436 38 438 43
rect 444 38 446 43
rect 460 38 462 43
rect 468 38 470 43
rect 484 38 486 43
<< ptransistor >>
rect 215 309 218 312
rect 231 309 234 312
rect 239 309 242 312
rect 255 309 258 312
rect 263 309 266 312
rect 279 309 282 312
rect 287 309 290 312
rect 303 309 306 312
rect 311 309 314 312
rect 327 309 330 312
rect 335 309 338 312
rect 351 309 354 312
rect 359 309 362 312
rect 375 309 378 312
rect 383 309 386 312
rect 399 309 402 312
rect 407 309 410 312
rect 423 309 426 312
rect 431 309 434 312
rect 447 309 450 312
rect 455 309 458 312
rect 471 309 474 312
rect 479 309 482 312
rect 14 275 17 278
rect 14 267 17 270
rect 14 251 17 254
rect 14 243 17 246
rect 14 227 17 230
rect 14 219 17 222
rect 14 203 17 206
rect 14 195 17 198
rect 14 179 17 182
rect 14 171 17 174
rect 14 155 17 158
rect 14 147 17 150
rect 14 131 17 134
rect 14 123 17 126
rect 14 107 17 110
rect 14 99 17 102
rect 14 83 17 86
rect 14 75 17 78
rect 14 59 17 62
rect 40 8 42 18
rect 56 8 58 18
rect 72 8 74 18
rect 88 8 90 18
rect 104 8 106 18
rect 120 8 122 18
rect 136 8 138 18
rect 152 8 154 18
rect 168 8 170 18
rect 184 8 186 18
rect 220 8 222 18
rect 228 8 230 18
rect 244 8 246 18
rect 252 8 254 18
rect 268 8 270 18
rect 276 8 278 18
rect 292 8 294 18
rect 300 8 302 18
rect 316 8 318 18
rect 324 8 326 18
rect 340 8 342 18
rect 348 8 350 18
rect 364 8 366 18
rect 372 8 374 18
rect 388 8 390 18
rect 396 8 398 18
rect 412 8 414 18
rect 420 8 422 18
rect 436 8 438 18
rect 444 8 446 18
rect 460 8 462 18
rect 468 8 470 18
rect 484 8 486 18
<< ndiffusion >>
rect 139 279 143 283
rect 155 279 159 283
rect 171 279 175 283
rect 43 183 47 187
rect 59 183 63 187
rect 43 179 48 183
rect 50 179 51 183
rect 55 179 56 183
rect 58 179 63 183
rect 43 171 48 175
rect 50 171 51 175
rect 55 171 56 175
rect 58 171 63 175
rect 43 167 47 171
rect 43 159 47 163
rect 39 155 40 159
rect 42 155 47 159
rect 39 147 40 151
rect 42 147 47 151
rect 43 143 47 147
rect 43 135 47 139
rect 39 131 40 135
rect 42 131 47 135
rect 59 167 63 171
rect 59 159 63 163
rect 55 155 56 159
rect 58 155 63 159
rect 55 147 56 151
rect 58 147 63 151
rect 59 143 63 147
rect 59 135 63 139
rect 55 131 56 135
rect 58 131 63 135
rect 43 123 48 127
rect 50 123 51 127
rect 55 123 56 127
rect 58 123 63 127
rect 43 119 47 123
rect 43 111 47 115
rect 59 119 63 123
rect 59 111 63 115
rect 43 107 48 111
rect 50 107 51 111
rect 55 107 56 111
rect 58 107 63 111
rect 35 42 40 43
rect 39 38 40 42
rect 42 42 47 43
rect 42 38 43 42
rect 51 42 56 43
rect 55 38 56 42
rect 58 42 63 43
rect 58 38 59 42
rect 75 183 79 187
rect 91 183 95 187
rect 75 179 80 183
rect 82 179 83 183
rect 87 179 88 183
rect 90 179 95 183
rect 71 171 72 175
rect 74 171 79 175
rect 75 167 79 171
rect 75 159 79 163
rect 71 155 72 159
rect 74 155 79 159
rect 71 147 72 151
rect 74 147 79 151
rect 75 143 79 147
rect 75 135 79 139
rect 71 131 72 135
rect 74 131 79 135
rect 87 171 88 175
rect 90 171 95 175
rect 91 167 95 171
rect 91 159 95 163
rect 87 155 88 159
rect 90 155 95 159
rect 107 183 111 187
rect 103 179 104 183
rect 106 179 111 183
rect 103 171 104 175
rect 106 171 111 175
rect 107 167 111 171
rect 107 159 111 163
rect 123 183 127 187
rect 119 179 120 183
rect 122 179 127 183
rect 119 171 120 175
rect 122 171 127 175
rect 123 167 127 171
rect 123 159 127 163
rect 107 155 112 159
rect 114 155 115 159
rect 119 155 120 159
rect 122 155 127 159
rect 91 147 96 151
rect 98 147 99 151
rect 103 147 104 151
rect 106 147 111 151
rect 91 143 95 147
rect 91 135 95 139
rect 87 131 88 135
rect 90 131 95 135
rect 75 123 80 127
rect 82 123 83 127
rect 87 123 88 127
rect 90 123 95 127
rect 75 119 79 123
rect 75 111 79 115
rect 71 107 72 111
rect 74 107 79 111
rect 67 42 72 43
rect 71 38 72 42
rect 74 42 79 43
rect 74 38 75 42
rect 91 119 95 123
rect 91 111 95 115
rect 87 107 88 111
rect 90 107 95 111
rect 83 42 88 43
rect 87 38 88 42
rect 90 42 95 43
rect 90 38 91 42
rect 107 143 111 147
rect 107 135 111 139
rect 103 131 104 135
rect 106 131 111 135
rect 103 123 104 127
rect 106 123 111 127
rect 107 119 111 123
rect 107 111 111 115
rect 103 107 104 111
rect 106 107 111 111
rect 99 42 104 43
rect 103 38 104 42
rect 106 42 111 43
rect 106 38 107 42
rect 119 147 120 151
rect 122 147 127 151
rect 123 143 127 147
rect 123 135 127 139
rect 119 131 120 135
rect 122 131 127 135
rect 119 123 120 127
rect 122 123 127 127
rect 123 119 127 123
rect 123 111 127 115
rect 119 107 120 111
rect 122 107 127 111
rect 115 42 120 43
rect 119 38 120 42
rect 122 42 127 43
rect 122 38 123 42
rect 139 275 144 279
rect 146 275 147 279
rect 139 267 144 271
rect 146 267 147 271
rect 139 263 143 267
rect 139 255 143 259
rect 155 275 160 279
rect 162 275 163 279
rect 167 275 168 279
rect 170 275 175 279
rect 187 279 191 283
rect 155 267 160 271
rect 162 267 163 271
rect 167 267 168 271
rect 170 267 175 271
rect 155 263 159 267
rect 155 255 159 259
rect 139 251 144 255
rect 146 251 147 255
rect 151 251 152 255
rect 154 251 159 255
rect 139 243 144 247
rect 146 243 147 247
rect 151 243 152 247
rect 154 243 159 247
rect 139 239 143 243
rect 139 231 143 235
rect 155 239 159 243
rect 155 231 159 235
rect 139 227 144 231
rect 146 227 147 231
rect 151 227 152 231
rect 154 227 159 231
rect 139 219 144 223
rect 146 219 147 223
rect 151 219 152 223
rect 154 219 159 223
rect 139 215 143 219
rect 139 207 143 211
rect 135 203 136 207
rect 138 203 143 207
rect 135 195 136 199
rect 138 195 143 199
rect 139 191 143 195
rect 139 183 143 187
rect 135 179 136 183
rect 138 179 143 183
rect 135 171 136 175
rect 138 171 143 175
rect 139 167 143 171
rect 139 159 143 163
rect 135 155 136 159
rect 138 155 143 159
rect 135 147 136 151
rect 138 147 143 151
rect 139 143 143 147
rect 139 135 143 139
rect 135 131 136 135
rect 138 131 143 135
rect 135 123 136 127
rect 138 123 143 127
rect 139 119 143 123
rect 139 111 143 115
rect 135 107 136 111
rect 138 107 143 111
rect 135 99 136 103
rect 138 99 143 103
rect 139 95 143 99
rect 139 87 143 91
rect 135 83 136 87
rect 138 83 143 87
rect 135 75 136 79
rect 138 75 143 79
rect 139 71 143 75
rect 139 63 143 67
rect 135 59 136 63
rect 138 59 143 63
rect 131 42 136 43
rect 135 38 136 42
rect 138 42 143 43
rect 138 38 139 42
rect 155 215 159 219
rect 155 207 159 211
rect 171 263 175 267
rect 171 255 175 259
rect 187 275 192 279
rect 194 275 195 279
rect 375 278 379 279
rect 375 275 379 276
rect 183 267 184 271
rect 186 267 191 271
rect 171 251 176 255
rect 178 251 179 255
rect 187 263 191 267
rect 187 255 191 259
rect 251 271 259 275
rect 255 270 259 271
rect 335 271 343 275
rect 371 271 379 275
rect 335 270 339 271
rect 255 267 259 268
rect 335 267 339 268
rect 187 251 192 255
rect 194 251 195 255
rect 231 254 235 255
rect 239 254 243 255
rect 351 254 355 255
rect 407 254 411 255
rect 231 251 235 252
rect 171 243 176 247
rect 178 243 179 247
rect 183 243 184 247
rect 186 243 191 247
rect 171 239 175 243
rect 171 231 175 235
rect 167 227 168 231
rect 170 227 175 231
rect 167 219 168 223
rect 170 219 175 223
rect 155 203 160 207
rect 162 203 163 207
rect 155 195 160 199
rect 162 195 163 199
rect 155 191 159 195
rect 155 183 159 187
rect 171 215 175 219
rect 171 207 175 211
rect 187 239 191 243
rect 187 231 191 235
rect 227 247 235 251
rect 239 251 243 252
rect 351 251 355 252
rect 407 251 411 252
rect 239 247 247 251
rect 347 247 355 251
rect 359 247 367 251
rect 371 247 379 251
rect 407 247 415 251
rect 359 246 363 247
rect 375 246 379 247
rect 359 243 363 244
rect 375 243 379 244
rect 187 227 192 231
rect 194 227 195 231
rect 215 230 219 231
rect 407 230 411 231
rect 447 230 451 231
rect 471 230 475 231
rect 215 227 219 228
rect 407 227 411 228
rect 447 227 451 228
rect 471 227 475 228
rect 183 219 184 223
rect 186 219 191 223
rect 171 203 176 207
rect 178 203 179 207
rect 187 215 191 219
rect 187 207 191 211
rect 215 223 223 227
rect 383 223 391 227
rect 407 223 415 227
rect 419 223 427 227
rect 443 223 451 227
rect 467 223 475 227
rect 383 222 387 223
rect 423 222 427 223
rect 383 219 387 220
rect 423 219 427 220
rect 187 203 192 207
rect 194 203 195 207
rect 375 206 379 207
rect 399 206 403 207
rect 375 203 379 204
rect 399 203 403 204
rect 171 195 176 199
rect 178 195 179 199
rect 183 195 184 199
rect 186 195 191 199
rect 171 191 175 195
rect 171 183 175 187
rect 155 179 160 183
rect 162 179 163 183
rect 167 179 168 183
rect 170 179 175 183
rect 155 171 160 175
rect 162 171 163 175
rect 167 171 168 175
rect 170 171 175 175
rect 155 167 159 171
rect 155 159 159 163
rect 171 167 175 171
rect 171 159 175 163
rect 155 155 160 159
rect 162 155 163 159
rect 167 155 168 159
rect 170 155 175 159
rect 155 147 160 151
rect 162 147 163 151
rect 167 147 168 151
rect 170 147 175 151
rect 155 143 159 147
rect 155 135 159 139
rect 171 143 175 147
rect 171 135 175 139
rect 155 131 160 135
rect 162 131 163 135
rect 167 131 168 135
rect 170 131 175 135
rect 155 123 160 127
rect 162 123 163 127
rect 167 123 168 127
rect 170 123 175 127
rect 155 119 159 123
rect 155 111 159 115
rect 171 119 175 123
rect 171 111 175 115
rect 155 107 160 111
rect 162 107 163 111
rect 167 107 168 111
rect 170 107 175 111
rect 151 99 152 103
rect 154 99 159 103
rect 155 95 159 99
rect 155 87 159 91
rect 151 83 152 87
rect 154 83 159 87
rect 151 75 152 79
rect 154 75 159 79
rect 155 71 159 75
rect 155 63 159 67
rect 151 59 152 63
rect 154 59 159 63
rect 147 42 152 43
rect 151 38 152 42
rect 154 42 159 43
rect 154 38 155 42
rect 187 191 191 195
rect 187 183 191 187
rect 371 199 379 203
rect 383 199 391 203
rect 395 199 403 203
rect 431 199 439 203
rect 455 199 463 203
rect 467 199 475 203
rect 383 198 387 199
rect 431 198 435 199
rect 455 198 459 199
rect 471 198 475 199
rect 479 199 487 203
rect 479 198 483 199
rect 383 195 387 196
rect 431 195 435 196
rect 455 195 459 196
rect 471 195 475 196
rect 479 195 483 196
rect 187 179 192 183
rect 194 179 195 183
rect 311 182 315 183
rect 407 182 411 183
rect 447 182 451 183
rect 311 179 315 180
rect 407 179 411 180
rect 447 179 451 180
rect 311 175 319 179
rect 407 175 415 179
rect 443 175 451 179
rect 455 175 463 179
rect 467 175 475 179
rect 187 171 192 175
rect 194 171 195 175
rect 311 174 315 175
rect 407 174 411 175
rect 455 174 459 175
rect 471 174 475 175
rect 311 171 315 172
rect 187 167 191 171
rect 187 159 191 163
rect 183 155 184 159
rect 186 155 191 159
rect 183 147 184 151
rect 186 147 191 151
rect 187 143 191 147
rect 187 135 191 139
rect 183 131 184 135
rect 186 131 191 135
rect 183 123 184 127
rect 186 123 191 127
rect 187 119 191 123
rect 187 111 191 115
rect 183 107 184 111
rect 186 107 191 111
rect 171 99 176 103
rect 178 99 179 103
rect 171 95 175 99
rect 171 87 175 91
rect 407 171 411 172
rect 455 171 459 172
rect 471 171 475 172
rect 311 158 315 159
rect 327 158 331 159
rect 447 158 451 159
rect 455 158 459 159
rect 311 155 315 156
rect 327 155 331 156
rect 447 155 451 156
rect 311 151 319 155
rect 323 151 331 155
rect 443 151 451 155
rect 455 155 459 156
rect 455 151 463 155
rect 467 151 475 155
rect 311 150 315 151
rect 327 150 331 151
rect 447 150 451 151
rect 471 150 475 151
rect 479 151 487 155
rect 479 150 483 151
rect 311 147 315 148
rect 327 147 331 148
rect 447 147 451 148
rect 471 147 475 148
rect 479 147 483 148
rect 311 134 315 135
rect 327 134 331 135
rect 447 134 451 135
rect 479 134 483 135
rect 311 131 315 132
rect 327 131 331 132
rect 447 131 451 132
rect 479 131 483 132
rect 311 127 319 131
rect 323 127 331 131
rect 443 127 451 131
rect 455 127 463 131
rect 479 127 487 131
rect 311 126 315 127
rect 327 126 331 127
rect 455 126 459 127
rect 479 126 483 127
rect 311 123 315 124
rect 327 123 331 124
rect 455 123 459 124
rect 479 123 483 124
rect 311 110 315 111
rect 327 110 331 111
rect 455 110 459 111
rect 479 110 483 111
rect 311 107 315 108
rect 327 107 331 108
rect 455 107 459 108
rect 479 107 483 108
rect 251 103 259 107
rect 187 99 192 103
rect 194 99 195 103
rect 255 102 259 103
rect 263 103 271 107
rect 311 103 319 107
rect 323 103 331 107
rect 263 102 267 103
rect 327 102 331 103
rect 431 103 439 107
rect 455 103 463 107
rect 479 103 487 107
rect 431 102 435 103
rect 455 102 459 103
rect 255 99 259 100
rect 187 95 191 99
rect 187 87 191 91
rect 171 83 176 87
rect 178 83 179 87
rect 183 83 184 87
rect 186 83 191 87
rect 167 75 168 79
rect 170 75 175 79
rect 171 71 175 75
rect 171 63 175 67
rect 167 59 168 63
rect 170 59 175 63
rect 163 42 168 43
rect 167 38 168 42
rect 170 42 175 43
rect 170 38 171 42
rect 263 99 267 100
rect 327 99 331 100
rect 431 99 435 100
rect 455 99 459 100
rect 255 86 259 87
rect 279 86 283 87
rect 327 86 331 87
rect 431 86 435 87
rect 471 86 475 87
rect 479 86 483 87
rect 255 83 259 84
rect 279 83 283 84
rect 327 83 331 84
rect 251 79 259 83
rect 275 79 283 83
rect 287 79 295 83
rect 323 79 331 83
rect 187 75 192 79
rect 194 75 195 79
rect 255 78 259 79
rect 287 78 291 79
rect 327 78 331 79
rect 431 83 435 84
rect 471 83 475 84
rect 431 79 439 83
rect 467 79 475 83
rect 479 83 483 84
rect 479 79 487 83
rect 431 78 435 79
rect 471 78 475 79
rect 255 75 259 76
rect 187 71 191 75
rect 187 63 191 67
rect 183 59 184 63
rect 186 59 191 63
rect 179 42 184 43
rect 183 38 184 42
rect 186 42 191 43
rect 186 38 187 42
rect 287 75 291 76
rect 327 75 331 76
rect 431 75 435 76
rect 471 75 475 76
rect 255 62 259 63
rect 303 62 307 63
rect 327 62 331 63
rect 431 62 435 63
rect 479 62 483 63
rect 255 59 259 60
rect 303 59 307 60
rect 327 59 331 60
rect 251 55 259 59
rect 299 55 307 59
rect 323 55 331 59
rect 431 59 435 60
rect 479 59 483 60
rect 431 55 439 59
rect 479 55 487 59
rect 215 42 220 43
rect 219 38 220 42
rect 222 42 228 43
rect 222 38 223 42
rect 227 38 228 42
rect 230 42 235 43
rect 230 38 231 42
rect 239 42 244 43
rect 243 38 244 42
rect 246 42 252 43
rect 246 38 247 42
rect 251 38 252 42
rect 254 42 259 43
rect 254 38 255 42
rect 263 42 268 43
rect 267 38 268 42
rect 270 42 276 43
rect 270 38 271 42
rect 275 38 276 42
rect 278 42 283 43
rect 278 38 279 42
rect 287 42 292 43
rect 291 38 292 42
rect 294 42 300 43
rect 294 38 295 42
rect 299 38 300 42
rect 302 42 307 43
rect 302 38 303 42
rect 311 42 316 43
rect 315 38 316 42
rect 318 42 324 43
rect 318 38 319 42
rect 323 38 324 42
rect 326 42 331 43
rect 326 38 327 42
rect 335 42 340 43
rect 339 38 340 42
rect 342 42 348 43
rect 342 38 343 42
rect 347 38 348 42
rect 350 42 355 43
rect 350 38 351 42
rect 359 42 364 43
rect 363 38 364 42
rect 366 42 372 43
rect 366 38 367 42
rect 371 38 372 42
rect 374 42 379 43
rect 374 38 375 42
rect 383 42 388 43
rect 387 38 388 42
rect 390 42 396 43
rect 390 38 391 42
rect 395 38 396 42
rect 398 42 403 43
rect 398 38 399 42
rect 407 42 412 43
rect 411 38 412 42
rect 414 42 420 43
rect 414 38 415 42
rect 419 38 420 42
rect 422 42 427 43
rect 422 38 423 42
rect 431 42 436 43
rect 435 38 436 42
rect 438 42 444 43
rect 438 38 439 42
rect 443 38 444 42
rect 446 42 451 43
rect 446 38 447 42
rect 455 42 460 43
rect 459 38 460 42
rect 462 42 468 43
rect 462 38 463 42
rect 467 38 468 42
rect 470 42 475 43
rect 470 38 471 42
rect 479 42 484 43
rect 483 38 484 42
rect 486 42 491 43
rect 486 38 487 42
<< pdiffusion >>
rect 215 312 218 314
rect 231 312 234 314
rect 239 312 242 314
rect 255 312 258 314
rect 263 312 266 314
rect 279 312 282 314
rect 287 312 290 314
rect 303 312 306 314
rect 311 312 314 314
rect 327 312 330 314
rect 335 312 338 314
rect 351 312 354 314
rect 359 312 362 314
rect 375 312 378 314
rect 383 312 386 314
rect 399 312 402 314
rect 407 312 410 314
rect 423 312 426 314
rect 431 312 434 314
rect 447 312 450 314
rect 455 312 458 314
rect 471 312 474 314
rect 479 312 482 314
rect 215 307 218 309
rect 231 307 234 309
rect 239 307 242 309
rect 255 307 258 309
rect 263 307 266 309
rect 279 307 282 309
rect 287 307 290 309
rect 303 307 306 309
rect 311 307 314 309
rect 327 307 330 309
rect 335 307 338 309
rect 351 307 354 309
rect 359 307 362 309
rect 375 307 378 309
rect 383 307 386 309
rect 399 307 402 309
rect 407 307 410 309
rect 423 307 426 309
rect 431 307 434 309
rect 447 307 450 309
rect 455 307 458 309
rect 471 307 474 309
rect 479 307 482 309
rect 12 275 14 278
rect 17 275 19 278
rect 12 267 14 270
rect 17 267 19 270
rect 12 251 14 254
rect 17 251 19 254
rect 12 243 14 246
rect 17 243 19 246
rect 12 227 14 230
rect 17 227 19 230
rect 12 219 14 222
rect 17 219 19 222
rect 12 203 14 206
rect 17 203 19 206
rect 12 195 14 198
rect 17 195 19 198
rect 12 179 14 182
rect 17 179 19 182
rect 12 171 14 174
rect 17 171 19 174
rect 12 155 14 158
rect 17 155 19 158
rect 12 147 14 150
rect 17 147 19 150
rect 12 131 14 134
rect 17 131 19 134
rect 12 123 14 126
rect 17 123 19 126
rect 12 107 14 110
rect 17 107 19 110
rect 12 99 14 102
rect 17 99 19 102
rect 12 83 14 86
rect 17 83 19 86
rect 12 75 14 78
rect 17 75 19 78
rect 12 59 14 62
rect 17 59 19 62
rect 35 17 40 18
rect 39 8 40 17
rect 42 17 47 18
rect 42 8 43 17
rect 51 17 56 18
rect 55 8 56 17
rect 58 17 63 18
rect 58 8 59 17
rect 67 17 72 18
rect 71 8 72 17
rect 74 17 79 18
rect 74 8 75 17
rect 83 17 88 18
rect 87 8 88 17
rect 90 17 95 18
rect 90 8 91 17
rect 99 17 104 18
rect 103 8 104 17
rect 106 17 111 18
rect 106 8 107 17
rect 115 17 120 18
rect 119 8 120 17
rect 122 17 127 18
rect 122 8 123 17
rect 131 17 136 18
rect 135 8 136 17
rect 138 17 143 18
rect 138 8 139 17
rect 147 17 152 18
rect 151 8 152 17
rect 154 17 159 18
rect 154 8 155 17
rect 163 17 168 18
rect 167 8 168 17
rect 170 17 175 18
rect 170 8 171 17
rect 179 17 184 18
rect 183 8 184 17
rect 186 17 191 18
rect 186 8 187 17
rect 215 17 220 18
rect 219 8 220 17
rect 222 17 228 18
rect 222 8 223 17
rect 227 8 228 17
rect 230 17 235 18
rect 230 8 231 17
rect 239 17 244 18
rect 243 8 244 17
rect 246 17 252 18
rect 246 8 247 17
rect 251 8 252 17
rect 254 17 259 18
rect 254 8 255 17
rect 263 17 268 18
rect 267 8 268 17
rect 270 17 276 18
rect 270 8 271 17
rect 275 8 276 17
rect 278 17 283 18
rect 278 8 279 17
rect 287 17 292 18
rect 291 8 292 17
rect 294 17 300 18
rect 294 8 295 17
rect 299 8 300 17
rect 302 17 307 18
rect 302 8 303 17
rect 311 17 316 18
rect 315 8 316 17
rect 318 17 324 18
rect 318 8 319 17
rect 323 8 324 17
rect 326 17 331 18
rect 326 8 327 17
rect 335 17 340 18
rect 339 8 340 17
rect 342 17 348 18
rect 342 8 343 17
rect 347 8 348 17
rect 350 17 355 18
rect 350 8 351 17
rect 359 17 364 18
rect 363 8 364 17
rect 366 17 372 18
rect 366 8 367 17
rect 371 8 372 17
rect 374 17 379 18
rect 374 8 375 17
rect 383 17 388 18
rect 387 8 388 17
rect 390 17 396 18
rect 390 8 391 17
rect 395 8 396 17
rect 398 17 403 18
rect 398 8 399 17
rect 407 17 412 18
rect 411 8 412 17
rect 414 17 420 18
rect 414 8 415 17
rect 419 8 420 17
rect 422 17 427 18
rect 422 8 423 17
rect 431 17 436 18
rect 435 8 436 17
rect 438 17 444 18
rect 438 8 439 17
rect 443 8 444 17
rect 446 17 451 18
rect 446 8 447 17
rect 455 17 460 18
rect 459 8 460 17
rect 462 17 468 18
rect 462 8 463 17
rect 467 8 468 17
rect 470 17 475 18
rect 470 8 471 17
rect 479 17 484 18
rect 483 8 484 17
rect 486 17 491 18
rect 486 8 487 17
<< ndcontact >>
rect 43 283 47 287
rect 59 283 63 287
rect 75 283 79 287
rect 91 283 95 287
rect 107 283 111 287
rect 123 283 127 287
rect 139 283 143 287
rect 155 283 159 287
rect 171 283 175 287
rect 187 283 191 287
rect 43 259 47 263
rect 43 235 47 239
rect 43 211 47 215
rect 43 187 47 191
rect 59 259 63 263
rect 59 235 63 239
rect 59 211 63 215
rect 59 187 63 191
rect 51 179 55 183
rect 51 171 55 175
rect 43 163 47 167
rect 35 155 39 159
rect 35 147 39 151
rect 43 139 47 143
rect 35 131 39 135
rect 59 163 63 167
rect 51 155 55 159
rect 51 147 55 151
rect 59 139 63 143
rect 51 131 55 135
rect 51 123 55 127
rect 43 115 47 119
rect 59 115 63 119
rect 51 107 55 111
rect 43 91 47 95
rect 43 67 47 71
rect 35 38 39 42
rect 43 38 47 42
rect 59 91 63 95
rect 59 67 63 71
rect 51 38 55 42
rect 59 38 63 42
rect 75 259 79 263
rect 75 235 79 239
rect 75 211 79 215
rect 75 187 79 191
rect 91 259 95 263
rect 91 235 95 239
rect 91 211 95 215
rect 91 187 95 191
rect 83 179 87 183
rect 67 171 71 175
rect 75 163 79 167
rect 67 155 71 159
rect 67 147 71 151
rect 75 139 79 143
rect 67 131 71 135
rect 83 171 87 175
rect 91 163 95 167
rect 83 155 87 159
rect 107 259 111 263
rect 107 235 111 239
rect 107 211 111 215
rect 107 187 111 191
rect 99 179 103 183
rect 99 171 103 175
rect 107 163 111 167
rect 123 259 127 263
rect 123 235 127 239
rect 123 211 127 215
rect 123 187 127 191
rect 115 179 119 183
rect 115 171 119 175
rect 123 163 127 167
rect 115 155 119 159
rect 99 147 103 151
rect 91 139 95 143
rect 83 131 87 135
rect 83 123 87 127
rect 75 115 79 119
rect 67 107 71 111
rect 75 91 79 95
rect 75 67 79 71
rect 67 38 71 42
rect 75 38 79 42
rect 91 115 95 119
rect 83 107 87 111
rect 91 91 95 95
rect 91 67 95 71
rect 83 38 87 42
rect 91 38 95 42
rect 107 139 111 143
rect 99 131 103 135
rect 99 123 103 127
rect 107 115 111 119
rect 99 107 103 111
rect 107 91 111 95
rect 107 67 111 71
rect 99 38 103 42
rect 107 38 111 42
rect 115 147 119 151
rect 123 139 127 143
rect 115 131 119 135
rect 115 123 119 127
rect 123 115 127 119
rect 115 107 119 111
rect 123 91 127 95
rect 123 67 127 71
rect 115 38 119 42
rect 123 38 127 42
rect 147 275 151 279
rect 147 267 151 271
rect 139 259 143 263
rect 163 275 167 279
rect 375 279 379 283
rect 163 267 167 271
rect 155 259 159 263
rect 147 251 151 255
rect 147 243 151 247
rect 139 235 143 239
rect 155 235 159 239
rect 147 227 151 231
rect 147 219 151 223
rect 139 211 143 215
rect 131 203 135 207
rect 131 195 135 199
rect 139 187 143 191
rect 131 179 135 183
rect 131 171 135 175
rect 139 163 143 167
rect 131 155 135 159
rect 131 147 135 151
rect 139 139 143 143
rect 131 131 135 135
rect 131 123 135 127
rect 139 115 143 119
rect 131 107 135 111
rect 131 99 135 103
rect 139 91 143 95
rect 131 83 135 87
rect 131 75 135 79
rect 139 67 143 71
rect 131 59 135 63
rect 131 38 135 42
rect 139 38 143 42
rect 155 211 159 215
rect 171 259 175 263
rect 195 275 199 279
rect 179 267 183 271
rect 179 251 183 255
rect 187 259 191 263
rect 247 271 251 275
rect 343 271 347 275
rect 367 271 371 275
rect 255 263 259 267
rect 335 263 339 267
rect 231 255 235 259
rect 195 251 199 255
rect 239 255 243 259
rect 351 255 355 259
rect 407 255 411 259
rect 179 243 183 247
rect 171 235 175 239
rect 163 227 167 231
rect 163 219 167 223
rect 163 203 167 207
rect 163 195 167 199
rect 155 187 159 191
rect 171 211 175 215
rect 187 235 191 239
rect 223 247 227 251
rect 247 247 251 251
rect 343 247 347 251
rect 367 247 371 251
rect 415 247 419 251
rect 359 239 363 243
rect 375 239 379 243
rect 215 231 219 235
rect 195 227 199 231
rect 407 231 411 235
rect 447 231 451 235
rect 471 231 475 235
rect 179 219 183 223
rect 179 203 183 207
rect 187 211 191 215
rect 223 223 227 227
rect 391 223 395 227
rect 415 223 419 227
rect 439 223 443 227
rect 463 223 467 227
rect 383 215 387 219
rect 423 215 427 219
rect 375 207 379 211
rect 195 203 199 207
rect 399 207 403 211
rect 179 195 183 199
rect 171 187 175 191
rect 163 179 167 183
rect 163 171 167 175
rect 155 163 159 167
rect 171 163 175 167
rect 163 155 167 159
rect 163 147 167 151
rect 155 139 159 143
rect 171 139 175 143
rect 163 131 167 135
rect 163 123 167 127
rect 155 115 159 119
rect 171 115 175 119
rect 163 107 167 111
rect 147 99 151 103
rect 155 91 159 95
rect 147 83 151 87
rect 147 75 151 79
rect 155 67 159 71
rect 147 59 151 63
rect 147 38 151 42
rect 155 38 159 42
rect 187 187 191 191
rect 367 199 371 203
rect 391 199 395 203
rect 439 199 443 203
rect 463 199 467 203
rect 487 199 491 203
rect 383 191 387 195
rect 431 191 435 195
rect 455 191 459 195
rect 471 191 475 195
rect 479 191 483 195
rect 311 183 315 187
rect 195 179 199 183
rect 407 183 411 187
rect 447 183 451 187
rect 319 175 323 179
rect 415 175 419 179
rect 439 175 443 179
rect 463 175 467 179
rect 195 171 199 175
rect 187 163 191 167
rect 179 155 183 159
rect 179 147 183 151
rect 187 139 191 143
rect 179 131 183 135
rect 179 123 183 127
rect 187 115 191 119
rect 179 107 183 111
rect 179 99 183 103
rect 171 91 175 95
rect 311 167 315 171
rect 407 167 411 171
rect 455 167 459 171
rect 471 167 475 171
rect 311 159 315 163
rect 327 159 331 163
rect 447 159 451 163
rect 455 159 459 163
rect 319 151 323 155
rect 439 151 443 155
rect 463 151 467 155
rect 487 151 491 155
rect 311 143 315 147
rect 327 143 331 147
rect 447 143 451 147
rect 471 143 475 147
rect 479 143 483 147
rect 311 135 315 139
rect 327 135 331 139
rect 447 135 451 139
rect 479 135 483 139
rect 319 127 323 131
rect 439 127 443 131
rect 463 127 467 131
rect 487 127 491 131
rect 311 119 315 123
rect 327 119 331 123
rect 455 119 459 123
rect 479 119 483 123
rect 311 111 315 115
rect 327 111 331 115
rect 455 111 459 115
rect 479 111 483 115
rect 247 103 251 107
rect 195 99 199 103
rect 271 103 275 107
rect 319 103 323 107
rect 439 103 443 107
rect 463 103 467 107
rect 487 103 491 107
rect 187 91 191 95
rect 179 83 183 87
rect 163 75 167 79
rect 171 67 175 71
rect 163 59 167 63
rect 163 38 167 42
rect 171 38 175 42
rect 255 95 259 99
rect 263 95 267 99
rect 327 95 331 99
rect 431 95 435 99
rect 455 95 459 99
rect 255 87 259 91
rect 279 87 283 91
rect 327 87 331 91
rect 431 87 435 91
rect 471 87 475 91
rect 479 87 483 91
rect 247 79 251 83
rect 271 79 275 83
rect 295 79 299 83
rect 319 79 323 83
rect 195 75 199 79
rect 439 79 443 83
rect 463 79 467 83
rect 487 79 491 83
rect 187 67 191 71
rect 179 59 183 63
rect 179 38 183 42
rect 187 38 191 42
rect 255 71 259 75
rect 287 71 291 75
rect 327 71 331 75
rect 431 71 435 75
rect 471 71 475 75
rect 255 63 259 67
rect 303 63 307 67
rect 327 63 331 67
rect 431 63 435 67
rect 479 63 483 67
rect 247 55 251 59
rect 295 55 299 59
rect 319 55 323 59
rect 439 55 443 59
rect 487 55 491 59
rect 215 38 219 42
rect 223 38 227 42
rect 231 38 235 42
rect 239 38 243 42
rect 247 38 251 42
rect 255 38 259 42
rect 263 38 267 42
rect 271 38 275 42
rect 279 38 283 42
rect 287 38 291 42
rect 295 38 299 42
rect 303 38 307 42
rect 311 38 315 42
rect 319 38 323 42
rect 327 38 331 42
rect 335 38 339 42
rect 343 38 347 42
rect 351 38 355 42
rect 359 38 363 42
rect 367 38 371 42
rect 375 38 379 42
rect 383 38 387 42
rect 391 38 395 42
rect 399 38 403 42
rect 407 38 411 42
rect 415 38 419 42
rect 423 38 427 42
rect 431 38 435 42
rect 439 38 443 42
rect 447 38 451 42
rect 455 38 459 42
rect 463 38 467 42
rect 471 38 475 42
rect 479 38 483 42
rect 487 38 491 42
<< pdcontact >>
rect 215 314 219 318
rect 231 314 235 318
rect 239 314 243 318
rect 255 314 259 318
rect 263 314 267 318
rect 279 314 283 318
rect 287 314 291 318
rect 303 314 307 318
rect 311 314 315 318
rect 327 314 331 318
rect 335 314 339 318
rect 351 314 355 318
rect 359 314 363 318
rect 375 314 379 318
rect 383 314 387 318
rect 399 314 403 318
rect 407 314 411 318
rect 423 314 427 318
rect 431 314 435 318
rect 447 314 451 318
rect 455 314 459 318
rect 471 314 475 318
rect 479 314 483 318
rect 215 303 219 307
rect 231 303 235 307
rect 239 303 243 307
rect 255 303 259 307
rect 263 303 267 307
rect 279 303 283 307
rect 287 303 291 307
rect 303 303 307 307
rect 311 303 315 307
rect 327 303 331 307
rect 335 303 339 307
rect 351 303 355 307
rect 359 303 363 307
rect 375 303 379 307
rect 383 303 387 307
rect 399 303 403 307
rect 407 303 411 307
rect 423 303 427 307
rect 431 303 435 307
rect 447 303 451 307
rect 455 303 459 307
rect 471 303 475 307
rect 479 303 483 307
rect 8 275 12 279
rect 19 275 23 279
rect 8 267 12 271
rect 19 267 23 271
rect 8 251 12 255
rect 19 251 23 255
rect 8 243 12 247
rect 19 243 23 247
rect 8 227 12 231
rect 19 227 23 231
rect 8 219 12 223
rect 19 219 23 223
rect 8 203 12 207
rect 19 203 23 207
rect 8 195 12 199
rect 19 195 23 199
rect 8 179 12 183
rect 19 179 23 183
rect 8 171 12 175
rect 19 171 23 175
rect 8 155 12 159
rect 19 155 23 159
rect 8 147 12 151
rect 19 147 23 151
rect 8 131 12 135
rect 19 131 23 135
rect 8 123 12 127
rect 19 123 23 127
rect 8 107 12 111
rect 19 107 23 111
rect 8 99 12 103
rect 19 99 23 103
rect 8 83 12 87
rect 19 83 23 87
rect 8 75 12 79
rect 19 75 23 79
rect 8 59 12 63
rect 19 59 23 63
rect 35 8 39 17
rect 43 8 47 17
rect 51 8 55 17
rect 59 8 63 17
rect 67 8 71 17
rect 75 8 79 17
rect 83 8 87 17
rect 91 8 95 17
rect 99 8 103 17
rect 107 8 111 17
rect 115 8 119 17
rect 123 8 127 17
rect 131 8 135 17
rect 139 8 143 17
rect 147 8 151 17
rect 155 8 159 17
rect 163 8 167 17
rect 171 8 175 17
rect 179 8 183 17
rect 187 8 191 17
rect 215 8 219 17
rect 223 8 227 17
rect 231 8 235 17
rect 239 8 243 17
rect 247 8 251 17
rect 255 8 259 17
rect 263 8 267 17
rect 271 8 275 17
rect 279 8 283 17
rect 287 8 291 17
rect 295 8 299 17
rect 303 8 307 17
rect 311 8 315 17
rect 319 8 323 17
rect 327 8 331 17
rect 335 8 339 17
rect 343 8 347 17
rect 351 8 355 17
rect 359 8 363 17
rect 367 8 371 17
rect 375 8 379 17
rect 383 8 387 17
rect 391 8 395 17
rect 399 8 403 17
rect 407 8 411 17
rect 415 8 419 17
rect 423 8 427 17
rect 431 8 435 17
rect 439 8 443 17
rect 447 8 451 17
rect 455 8 459 17
rect 463 8 467 17
rect 471 8 475 17
rect 479 8 483 17
rect 487 8 491 17
<< psubstratepcontact >>
rect 35 283 39 287
rect 51 283 55 287
rect 67 283 71 287
rect 83 283 87 287
rect 99 283 103 287
rect 115 283 119 287
rect 131 283 135 287
rect 147 283 151 287
rect 163 283 167 287
rect 179 283 183 287
rect 195 283 199 287
rect 223 283 227 287
rect 247 283 251 287
rect 271 283 275 287
rect 295 283 299 287
rect 319 283 323 287
rect 343 283 347 287
rect 367 283 371 287
rect 391 283 395 287
rect 415 283 419 287
rect 439 283 443 287
rect 463 283 467 287
rect 487 283 491 287
rect 35 259 39 263
rect 35 235 39 239
rect 35 211 39 215
rect 35 187 39 191
rect 35 163 39 167
rect 51 259 55 263
rect 51 235 55 239
rect 51 211 55 215
rect 51 187 55 191
rect 35 139 39 143
rect 35 115 39 119
rect 35 91 39 95
rect 35 67 39 71
rect 35 49 39 53
rect 51 163 55 167
rect 51 139 55 143
rect 51 115 55 119
rect 51 91 55 95
rect 51 67 55 71
rect 51 49 55 53
rect 67 259 71 263
rect 67 235 71 239
rect 67 211 71 215
rect 67 187 71 191
rect 83 259 87 263
rect 83 235 87 239
rect 83 211 87 215
rect 83 187 87 191
rect 67 163 71 167
rect 67 139 71 143
rect 67 115 71 119
rect 83 163 87 167
rect 83 139 87 143
rect 99 259 103 263
rect 99 235 103 239
rect 99 211 103 215
rect 99 187 103 191
rect 99 163 103 167
rect 115 259 119 263
rect 115 235 119 239
rect 115 211 119 215
rect 115 187 119 191
rect 115 163 119 167
rect 67 91 71 95
rect 67 67 71 71
rect 67 49 71 53
rect 83 115 87 119
rect 83 91 87 95
rect 83 67 87 71
rect 83 49 87 53
rect 99 139 103 143
rect 99 115 103 119
rect 99 91 103 95
rect 99 67 103 71
rect 99 49 103 53
rect 115 139 119 143
rect 115 115 119 119
rect 115 91 119 95
rect 115 67 119 71
rect 115 49 119 53
rect 131 259 135 263
rect 131 235 135 239
rect 131 211 135 215
rect 147 259 151 263
rect 147 235 151 239
rect 131 187 135 191
rect 131 163 135 167
rect 131 139 135 143
rect 131 115 135 119
rect 131 91 135 95
rect 131 67 135 71
rect 131 49 135 53
rect 147 211 151 215
rect 147 187 151 191
rect 147 163 151 167
rect 147 139 151 143
rect 147 115 151 119
rect 163 259 167 263
rect 163 235 167 239
rect 179 259 183 263
rect 195 259 199 263
rect 223 259 227 263
rect 247 259 251 263
rect 271 259 275 263
rect 295 259 299 263
rect 319 259 323 263
rect 343 259 347 263
rect 367 259 371 263
rect 391 259 395 263
rect 415 259 419 263
rect 439 259 443 263
rect 463 259 467 263
rect 487 259 491 263
rect 163 211 167 215
rect 163 187 167 191
rect 179 235 183 239
rect 195 235 199 239
rect 223 235 227 239
rect 247 235 251 239
rect 271 235 275 239
rect 295 235 299 239
rect 319 235 323 239
rect 343 235 347 239
rect 367 235 371 239
rect 391 235 395 239
rect 415 235 419 239
rect 439 235 443 239
rect 463 235 467 239
rect 487 235 491 239
rect 179 211 183 215
rect 195 211 199 215
rect 223 211 227 215
rect 247 211 251 215
rect 271 211 275 215
rect 295 211 299 215
rect 319 211 323 215
rect 343 211 347 215
rect 367 211 371 215
rect 391 211 395 215
rect 415 211 419 215
rect 439 211 443 215
rect 463 211 467 215
rect 487 211 491 215
rect 163 163 167 167
rect 163 139 167 143
rect 163 115 167 119
rect 147 91 151 95
rect 147 67 151 71
rect 147 49 151 53
rect 163 91 167 95
rect 179 187 183 191
rect 179 163 183 167
rect 195 187 199 191
rect 223 187 227 191
rect 247 187 251 191
rect 271 187 275 191
rect 295 187 299 191
rect 319 187 323 191
rect 343 187 347 191
rect 367 187 371 191
rect 391 187 395 191
rect 415 187 419 191
rect 439 187 443 191
rect 463 187 467 191
rect 487 187 491 191
rect 179 139 183 143
rect 179 115 183 119
rect 179 91 183 95
rect 195 163 199 167
rect 223 163 227 167
rect 247 163 251 167
rect 271 163 275 167
rect 295 163 299 167
rect 319 163 323 167
rect 343 163 347 167
rect 367 163 371 167
rect 391 163 395 167
rect 415 163 419 167
rect 439 163 443 167
rect 463 163 467 167
rect 487 163 491 167
rect 195 139 199 143
rect 223 139 227 143
rect 247 139 251 143
rect 271 139 275 143
rect 295 139 299 143
rect 319 139 323 143
rect 343 139 347 143
rect 367 139 371 143
rect 391 139 395 143
rect 415 139 419 143
rect 439 139 443 143
rect 463 139 467 143
rect 487 139 491 143
rect 195 115 199 119
rect 223 115 227 119
rect 247 115 251 119
rect 271 115 275 119
rect 295 115 299 119
rect 319 115 323 119
rect 343 115 347 119
rect 367 115 371 119
rect 391 115 395 119
rect 415 115 419 119
rect 439 115 443 119
rect 463 115 467 119
rect 487 115 491 119
rect 163 67 167 71
rect 163 49 167 53
rect 179 67 183 71
rect 195 91 199 95
rect 223 91 227 95
rect 247 91 251 95
rect 271 91 275 95
rect 295 91 299 95
rect 319 91 323 95
rect 343 91 347 95
rect 367 91 371 95
rect 391 91 395 95
rect 415 91 419 95
rect 439 91 443 95
rect 463 91 467 95
rect 487 91 491 95
rect 179 49 183 53
rect 195 67 199 71
rect 223 67 227 71
rect 247 67 251 71
rect 271 67 275 71
rect 295 67 299 71
rect 319 67 323 71
rect 343 67 347 71
rect 367 67 371 71
rect 391 67 395 71
rect 415 67 419 71
rect 439 67 443 71
rect 463 67 467 71
rect 487 67 491 71
<< nsubstratencontact >>
rect 215 322 219 326
rect 223 322 227 326
rect 231 322 235 326
rect 239 322 243 326
rect 247 322 251 326
rect 255 322 259 326
rect 263 322 267 326
rect 271 322 275 326
rect 279 322 283 326
rect 287 322 291 326
rect 295 322 299 326
rect 303 322 307 326
rect 311 322 315 326
rect 319 322 323 326
rect 327 322 331 326
rect 335 322 339 326
rect 343 322 347 326
rect 351 322 355 326
rect 359 322 363 326
rect 367 322 371 326
rect 375 322 379 326
rect 383 322 387 326
rect 391 322 395 326
rect 399 322 403 326
rect 407 322 411 326
rect 415 322 419 326
rect 423 322 427 326
rect 431 322 435 326
rect 439 322 443 326
rect 447 322 451 326
rect 455 322 459 326
rect 463 322 467 326
rect 471 322 475 326
rect 479 322 483 326
rect 487 322 491 326
rect 0 275 4 279
rect 0 267 4 271
rect 0 259 4 263
rect 0 251 4 255
rect 0 243 4 247
rect 0 235 4 239
rect 0 227 4 231
rect 0 219 4 223
rect 0 211 4 215
rect 0 203 4 207
rect 0 195 4 199
rect 0 187 4 191
rect 0 179 4 183
rect 0 171 4 175
rect 0 163 4 167
rect 0 155 4 159
rect 0 147 4 151
rect 0 139 4 143
rect 0 131 4 135
rect 0 123 4 127
rect 0 115 4 119
rect 0 107 4 111
rect 0 99 4 103
rect 0 91 4 95
rect 0 83 4 87
rect 0 75 4 79
rect 0 67 4 71
rect 0 59 4 63
rect 35 -2 39 2
rect 43 -2 47 2
rect 51 -2 55 2
rect 59 -2 63 2
rect 67 -2 71 2
rect 75 -2 79 2
rect 83 -2 87 2
rect 91 -2 95 2
rect 99 -2 103 2
rect 107 -2 111 2
rect 115 -2 119 2
rect 123 -2 127 2
rect 131 -2 135 2
rect 139 -2 143 2
rect 147 -2 151 2
rect 155 -2 159 2
rect 163 -2 167 2
rect 171 -2 175 2
rect 179 -2 183 2
rect 187 -2 191 2
rect 215 -2 219 2
rect 223 -2 227 2
rect 231 -2 235 2
rect 239 -2 243 2
rect 247 -2 251 2
rect 255 -2 259 2
rect 263 -2 267 2
rect 271 -2 275 2
rect 279 -2 283 2
rect 287 -2 291 2
rect 295 -2 299 2
rect 303 -2 307 2
rect 311 -2 315 2
rect 319 -2 323 2
rect 327 -2 331 2
rect 335 -2 339 2
rect 343 -2 347 2
rect 351 -2 355 2
rect 359 -2 363 2
rect 367 -2 371 2
rect 375 -2 379 2
rect 383 -2 387 2
rect 391 -2 395 2
rect 399 -2 403 2
rect 407 -2 411 2
rect 415 -2 419 2
rect 423 -2 427 2
rect 431 -2 435 2
rect 439 -2 443 2
rect 447 -2 451 2
rect 455 -2 459 2
rect 463 -2 467 2
rect 471 -2 475 2
rect 479 -2 483 2
rect 487 -2 491 2
<< polysilicon >>
rect 213 309 215 312
rect 218 309 223 312
rect 227 309 231 312
rect 234 309 239 312
rect 242 309 247 312
rect 251 309 255 312
rect 258 309 263 312
rect 266 309 271 312
rect 275 309 279 312
rect 282 309 287 312
rect 290 309 295 312
rect 299 309 303 312
rect 306 309 311 312
rect 314 309 319 312
rect 323 309 327 312
rect 330 309 335 312
rect 338 309 343 312
rect 347 309 351 312
rect 354 309 359 312
rect 362 309 367 312
rect 371 309 375 312
rect 378 309 383 312
rect 386 309 391 312
rect 395 309 399 312
rect 402 309 407 312
rect 410 309 415 312
rect 419 309 423 312
rect 426 309 431 312
rect 434 309 439 312
rect 443 309 447 312
rect 450 309 455 312
rect 458 309 463 312
rect 467 309 471 312
rect 474 309 479 312
rect 482 309 487 312
rect 14 278 17 283
rect 144 279 146 281
rect 160 279 162 281
rect 168 279 170 281
rect 14 270 17 275
rect 14 263 17 267
rect 14 254 17 259
rect 14 246 17 251
rect 14 239 17 243
rect 14 230 17 235
rect 14 222 17 227
rect 14 215 17 219
rect 14 206 17 211
rect 14 198 17 203
rect 14 191 17 195
rect 14 182 17 187
rect 14 174 17 179
rect 14 167 17 171
rect 14 158 17 163
rect 40 159 42 278
rect 48 183 50 278
rect 56 183 58 278
rect 48 175 50 179
rect 56 175 58 179
rect 14 150 17 155
rect 40 151 42 155
rect 14 143 17 147
rect 14 134 17 139
rect 40 135 42 147
rect 14 126 17 131
rect 14 119 17 123
rect 14 110 17 115
rect 14 102 17 107
rect 14 95 17 99
rect 14 86 17 91
rect 14 78 17 83
rect 14 71 17 75
rect 14 62 17 67
rect 14 57 17 59
rect 40 43 42 131
rect 48 127 50 171
rect 56 159 58 171
rect 56 151 58 155
rect 56 135 58 147
rect 56 127 58 131
rect 48 111 50 123
rect 56 111 58 123
rect 40 28 42 38
rect 48 34 50 107
rect 56 43 58 107
rect 56 28 58 38
rect 64 34 66 278
rect 72 175 74 278
rect 80 183 82 278
rect 88 183 90 278
rect 72 159 74 171
rect 72 151 74 155
rect 72 135 74 147
rect 72 111 74 131
rect 80 127 82 179
rect 88 175 90 179
rect 88 159 90 171
rect 88 135 90 155
rect 96 151 98 278
rect 104 183 106 278
rect 104 175 106 179
rect 104 151 106 171
rect 112 159 114 278
rect 120 183 122 278
rect 120 175 122 179
rect 120 159 122 171
rect 88 127 90 131
rect 72 43 74 107
rect 72 28 74 38
rect 80 34 82 123
rect 88 111 90 123
rect 88 43 90 107
rect 88 28 90 38
rect 96 34 98 147
rect 104 135 106 147
rect 104 127 106 131
rect 104 111 106 123
rect 104 43 106 107
rect 104 28 106 38
rect 112 34 114 155
rect 120 151 122 155
rect 120 135 122 147
rect 120 127 122 131
rect 120 111 122 123
rect 120 43 122 107
rect 120 28 122 38
rect 128 34 130 278
rect 136 207 138 278
rect 144 271 146 275
rect 144 255 146 267
rect 152 255 154 278
rect 192 279 194 281
rect 160 271 162 275
rect 168 271 170 275
rect 144 247 146 251
rect 152 247 154 251
rect 144 231 146 243
rect 152 231 154 243
rect 144 223 146 227
rect 152 223 154 227
rect 136 199 138 203
rect 136 183 138 195
rect 136 175 138 179
rect 136 159 138 171
rect 136 151 138 155
rect 136 135 138 147
rect 136 127 138 131
rect 136 111 138 123
rect 136 103 138 107
rect 136 87 138 99
rect 136 79 138 83
rect 136 63 138 75
rect 136 43 138 59
rect 136 28 138 38
rect 144 34 146 219
rect 152 103 154 219
rect 160 207 162 267
rect 168 231 170 267
rect 176 255 178 278
rect 184 271 186 278
rect 209 276 375 278
rect 379 276 482 278
rect 176 247 178 251
rect 184 247 186 267
rect 192 255 194 275
rect 209 268 255 270
rect 259 268 335 270
rect 339 268 482 270
rect 209 252 231 254
rect 235 252 239 254
rect 243 252 351 254
rect 355 252 407 254
rect 411 252 482 254
rect 168 223 170 227
rect 160 199 162 203
rect 160 183 162 195
rect 168 183 170 219
rect 176 207 178 243
rect 184 223 186 243
rect 192 231 194 251
rect 209 244 359 246
rect 363 244 375 246
rect 379 244 482 246
rect 209 228 215 230
rect 219 228 407 230
rect 411 228 447 230
rect 451 228 471 230
rect 475 228 482 230
rect 176 199 178 203
rect 184 199 186 219
rect 192 207 194 227
rect 209 220 383 222
rect 387 220 423 222
rect 427 220 482 222
rect 209 204 375 206
rect 379 204 399 206
rect 403 204 482 206
rect 160 175 162 179
rect 168 175 170 179
rect 160 159 162 171
rect 168 159 170 171
rect 160 151 162 155
rect 168 151 170 155
rect 160 135 162 147
rect 168 135 170 147
rect 160 127 162 131
rect 168 127 170 131
rect 160 111 162 123
rect 168 111 170 123
rect 152 87 154 99
rect 152 79 154 83
rect 152 63 154 75
rect 152 43 154 59
rect 152 28 154 38
rect 160 34 162 107
rect 168 79 170 107
rect 176 103 178 195
rect 184 159 186 195
rect 192 183 194 203
rect 209 196 383 198
rect 387 196 431 198
rect 435 196 455 198
rect 459 196 471 198
rect 475 196 479 198
rect 483 196 485 198
rect 209 180 311 182
rect 315 180 407 182
rect 411 180 447 182
rect 451 180 482 182
rect 192 175 194 179
rect 209 172 311 174
rect 315 172 407 174
rect 411 172 455 174
rect 459 172 471 174
rect 475 172 482 174
rect 184 151 186 155
rect 184 135 186 147
rect 184 127 186 131
rect 184 111 186 123
rect 176 87 178 99
rect 184 87 186 107
rect 192 103 194 171
rect 209 156 311 158
rect 315 156 327 158
rect 331 156 447 158
rect 451 156 455 158
rect 459 156 482 158
rect 209 148 311 150
rect 315 148 327 150
rect 331 148 447 150
rect 451 148 471 150
rect 475 148 479 150
rect 483 148 485 150
rect 209 132 311 134
rect 315 132 327 134
rect 331 132 447 134
rect 451 132 479 134
rect 483 132 485 134
rect 209 124 311 126
rect 315 124 327 126
rect 331 124 455 126
rect 459 124 479 126
rect 483 124 485 126
rect 209 108 311 110
rect 315 108 327 110
rect 331 108 455 110
rect 459 108 479 110
rect 483 108 485 110
rect 209 100 255 102
rect 259 100 263 102
rect 267 100 327 102
rect 331 100 431 102
rect 435 100 455 102
rect 459 100 482 102
rect 168 63 170 75
rect 168 43 170 59
rect 168 28 170 38
rect 176 34 178 83
rect 184 63 186 83
rect 192 79 194 99
rect 209 84 255 86
rect 259 84 279 86
rect 283 84 327 86
rect 331 84 431 86
rect 435 84 471 86
rect 475 84 479 86
rect 483 84 485 86
rect 209 76 255 78
rect 259 76 287 78
rect 291 76 327 78
rect 331 76 431 78
rect 435 76 471 78
rect 475 76 482 78
rect 184 43 186 59
rect 184 28 186 38
rect 192 34 194 75
rect 209 60 255 62
rect 259 60 303 62
rect 307 60 327 62
rect 331 60 431 62
rect 435 60 479 62
rect 483 60 485 62
rect 220 43 222 52
rect 228 43 230 52
rect 244 43 246 52
rect 252 43 254 52
rect 268 43 270 52
rect 276 43 278 52
rect 292 43 294 52
rect 300 43 302 52
rect 316 43 318 52
rect 324 43 326 52
rect 340 43 342 52
rect 348 43 350 52
rect 364 43 366 52
rect 372 43 374 52
rect 388 43 390 52
rect 396 43 398 52
rect 412 43 414 52
rect 420 43 422 52
rect 436 43 438 52
rect 444 43 446 52
rect 460 43 462 52
rect 468 43 470 52
rect 484 43 486 52
rect 37 26 42 28
rect 54 26 58 28
rect 70 26 74 28
rect 86 26 90 28
rect 102 26 106 28
rect 118 26 122 28
rect 134 26 138 28
rect 150 26 154 28
rect 166 26 170 28
rect 182 26 186 28
rect 83 22 84 26
rect 37 20 42 22
rect 54 20 58 22
rect 69 20 74 22
rect 85 20 90 22
rect 101 20 106 22
rect 117 20 122 22
rect 133 20 138 22
rect 149 20 154 22
rect 165 20 170 22
rect 181 20 186 22
rect 40 18 42 20
rect 56 18 58 20
rect 72 18 74 20
rect 88 18 90 20
rect 104 18 106 20
rect 120 18 122 20
rect 136 18 138 20
rect 152 18 154 20
rect 168 18 170 20
rect 184 18 186 20
rect 220 18 222 38
rect 228 18 230 38
rect 244 18 246 38
rect 252 18 254 38
rect 268 18 270 38
rect 276 18 278 38
rect 292 18 294 38
rect 300 18 302 38
rect 316 18 318 38
rect 324 18 326 38
rect 340 18 342 38
rect 348 18 350 38
rect 364 18 366 38
rect 372 18 374 38
rect 388 18 390 38
rect 396 18 398 38
rect 412 18 414 38
rect 420 18 422 38
rect 436 18 438 38
rect 444 18 446 38
rect 460 18 462 38
rect 468 18 470 38
rect 484 18 486 38
rect 40 6 42 8
rect 56 6 58 8
rect 72 6 74 8
rect 88 6 90 8
rect 104 6 106 8
rect 120 6 122 8
rect 136 6 138 8
rect 152 6 154 8
rect 168 6 170 8
rect 184 6 186 8
rect 220 6 222 8
rect 228 6 230 8
rect 244 6 246 8
rect 252 6 254 8
rect 268 6 270 8
rect 276 6 278 8
rect 292 6 294 8
rect 300 6 302 8
rect 316 6 318 8
rect 324 6 326 8
rect 340 6 342 8
rect 348 6 350 8
rect 364 6 366 8
rect 372 6 374 8
rect 388 6 390 8
rect 396 6 398 8
rect 412 6 414 8
rect 420 6 422 8
rect 436 6 438 8
rect 444 6 446 8
rect 460 6 462 8
rect 468 6 470 8
rect 484 6 486 8
<< polycontact >>
rect 223 308 227 312
rect 247 308 251 312
rect 271 308 275 312
rect 295 308 299 312
rect 319 308 323 312
rect 343 308 347 312
rect 367 308 371 312
rect 391 308 395 312
rect 415 308 419 312
rect 439 308 443 312
rect 463 308 467 312
rect 487 308 491 312
rect 13 283 17 287
rect 13 259 17 263
rect 13 235 17 239
rect 13 211 17 215
rect 13 187 17 191
rect 13 163 17 167
rect 13 139 17 143
rect 13 115 17 119
rect 13 91 17 95
rect 13 67 17 71
rect 46 30 50 34
rect 62 30 66 34
rect 78 30 82 34
rect 94 30 98 34
rect 110 30 114 34
rect 126 30 130 34
rect 205 275 209 279
rect 205 267 209 271
rect 205 251 209 255
rect 205 243 209 247
rect 205 227 209 231
rect 205 219 209 223
rect 205 203 209 207
rect 142 30 146 34
rect 205 195 209 199
rect 205 179 209 183
rect 205 171 209 175
rect 205 155 209 159
rect 205 147 209 151
rect 205 131 209 135
rect 205 123 209 127
rect 205 107 209 111
rect 205 99 209 103
rect 158 30 162 34
rect 205 83 209 87
rect 205 75 209 79
rect 174 30 178 34
rect 205 59 209 63
rect 216 49 220 53
rect 230 49 234 53
rect 240 49 244 53
rect 254 49 258 53
rect 264 49 268 53
rect 278 49 282 53
rect 288 49 292 53
rect 302 49 306 53
rect 312 49 316 53
rect 326 49 330 53
rect 336 49 340 53
rect 350 49 354 53
rect 360 49 364 53
rect 374 49 378 53
rect 384 49 388 53
rect 398 49 402 53
rect 408 49 412 53
rect 422 49 426 53
rect 432 49 436 53
rect 446 49 450 53
rect 456 49 460 53
rect 470 49 474 53
rect 480 49 484 53
rect 190 30 194 34
rect 35 22 39 26
rect 51 22 56 26
rect 67 22 72 26
rect 84 22 88 26
rect 100 22 104 26
rect 116 22 120 26
rect 132 22 136 26
rect 148 22 152 26
rect 164 22 168 26
rect 180 22 184 26
<< metal1 >>
rect 203 338 493 340
rect 203 334 205 338
rect 209 334 223 338
rect 227 334 247 338
rect 251 334 271 338
rect 275 334 295 338
rect 299 334 319 338
rect 323 334 343 338
rect 347 334 367 338
rect 371 334 391 338
rect 395 334 415 338
rect 419 334 439 338
rect 443 334 463 338
rect 467 334 487 338
rect 491 334 493 338
rect 203 332 493 334
rect -2 326 493 328
rect -2 322 215 326
rect 219 322 223 326
rect 227 322 231 326
rect 235 322 239 326
rect 243 322 247 326
rect 251 322 255 326
rect 259 322 263 326
rect 267 322 271 326
rect 275 322 279 326
rect 283 322 287 326
rect 291 322 295 326
rect 299 322 303 326
rect 307 322 311 326
rect 315 322 319 326
rect 323 322 327 326
rect 331 322 335 326
rect 339 322 343 326
rect 347 322 351 326
rect 355 322 359 326
rect 363 322 367 326
rect 371 322 375 326
rect 379 322 383 326
rect 387 322 391 326
rect 395 322 399 326
rect 403 322 407 326
rect 411 322 415 326
rect 419 322 423 326
rect 427 322 431 326
rect 435 322 439 326
rect 443 322 447 326
rect 451 322 455 326
rect 459 322 463 326
rect 467 322 471 326
rect 475 322 479 326
rect 483 322 487 326
rect 491 322 493 326
rect -2 320 493 322
rect -2 279 6 320
rect 215 318 219 320
rect 231 318 235 320
rect 239 318 243 320
rect 255 318 259 320
rect 263 318 267 320
rect 279 318 283 320
rect 287 318 291 320
rect 303 318 307 320
rect 311 318 315 320
rect 327 318 331 320
rect 335 318 339 320
rect 351 318 355 320
rect 359 318 363 320
rect 375 318 379 320
rect 383 318 387 320
rect 399 318 403 320
rect 407 318 411 320
rect 423 318 427 320
rect 431 318 435 320
rect 447 318 451 320
rect 455 318 459 320
rect 471 318 475 320
rect 479 318 483 320
rect 17 283 35 287
rect 39 283 43 287
rect 47 283 51 287
rect 55 283 59 287
rect 63 283 67 287
rect 71 283 75 287
rect 79 283 83 287
rect 87 283 91 287
rect 95 283 99 287
rect 103 283 107 287
rect 111 283 115 287
rect 119 283 123 287
rect 127 283 131 287
rect 135 283 139 287
rect 143 283 147 287
rect 151 283 155 287
rect 159 283 163 287
rect 167 283 171 287
rect 175 283 179 287
rect 183 283 187 287
rect 191 283 195 287
rect 199 283 205 287
rect -2 275 0 279
rect 4 275 8 279
rect 23 275 147 279
rect 151 275 163 279
rect 167 275 195 279
rect 199 275 205 279
rect -2 271 6 275
rect -2 267 0 271
rect 4 267 8 271
rect 23 267 147 271
rect 151 267 163 271
rect 167 267 179 271
rect 183 267 205 271
rect -2 263 6 267
rect -2 259 0 263
rect 4 259 6 263
rect 17 259 35 263
rect 39 259 43 263
rect 47 259 51 263
rect 55 259 59 263
rect 63 259 67 263
rect 71 259 75 263
rect 79 259 83 263
rect 87 259 91 263
rect 95 259 99 263
rect 103 259 107 263
rect 111 259 115 263
rect 119 259 123 263
rect 127 259 131 263
rect 135 259 139 263
rect 143 259 147 263
rect 151 259 155 263
rect 159 259 163 263
rect 167 259 171 263
rect 175 259 179 263
rect 183 259 187 263
rect 191 259 195 263
rect 199 259 205 263
rect -2 255 6 259
rect -2 251 0 255
rect 4 251 8 255
rect 23 251 147 255
rect 151 251 179 255
rect 183 251 195 255
rect 199 251 205 255
rect -2 247 6 251
rect -2 243 0 247
rect 4 243 8 247
rect 23 243 147 247
rect 151 243 179 247
rect 183 243 205 247
rect -2 239 6 243
rect -2 235 0 239
rect 4 235 6 239
rect 17 235 35 239
rect 39 235 43 239
rect 47 235 51 239
rect 55 235 59 239
rect 63 235 67 239
rect 71 235 75 239
rect 79 235 83 239
rect 87 235 91 239
rect 95 235 99 239
rect 103 235 107 239
rect 111 235 115 239
rect 119 235 123 239
rect 127 235 131 239
rect 135 235 139 239
rect 143 235 147 239
rect 151 235 155 239
rect 159 235 163 239
rect 167 235 171 239
rect 175 235 179 239
rect 183 235 187 239
rect 191 235 195 239
rect 199 235 205 239
rect 215 235 219 303
rect -2 231 6 235
rect -2 227 0 231
rect 4 227 8 231
rect 23 227 147 231
rect 151 227 163 231
rect 167 227 195 231
rect 199 227 205 231
rect -2 223 6 227
rect -2 219 0 223
rect 4 219 8 223
rect 23 219 147 223
rect 151 219 163 223
rect 167 219 179 223
rect 183 219 205 223
rect -2 215 6 219
rect -2 211 0 215
rect 4 211 6 215
rect 17 211 35 215
rect 39 211 43 215
rect 47 211 51 215
rect 55 211 59 215
rect 63 211 67 215
rect 71 211 75 215
rect 79 211 83 215
rect 87 211 91 215
rect 95 211 99 215
rect 103 211 107 215
rect 111 211 115 215
rect 119 211 123 215
rect 127 211 131 215
rect 135 211 139 215
rect 143 211 147 215
rect 151 211 155 215
rect 159 211 163 215
rect 167 211 171 215
rect 175 211 179 215
rect 183 211 187 215
rect 191 211 195 215
rect 199 211 205 215
rect -2 207 6 211
rect -2 203 0 207
rect 4 203 8 207
rect 23 203 131 207
rect 135 203 163 207
rect 167 203 179 207
rect 183 203 195 207
rect 199 203 205 207
rect -2 199 6 203
rect -2 195 0 199
rect 4 195 8 199
rect 23 195 131 199
rect 135 195 163 199
rect 167 195 179 199
rect 183 195 205 199
rect -2 191 6 195
rect -2 187 0 191
rect 4 187 6 191
rect 17 187 35 191
rect 39 187 43 191
rect 47 187 51 191
rect 55 187 59 191
rect 63 187 67 191
rect 71 187 75 191
rect 79 187 83 191
rect 87 187 91 191
rect 95 187 99 191
rect 103 187 107 191
rect 111 187 115 191
rect 119 187 123 191
rect 127 187 131 191
rect 135 187 139 191
rect 143 187 147 191
rect 151 187 155 191
rect 159 187 163 191
rect 167 187 171 191
rect 175 187 179 191
rect 183 187 187 191
rect 191 187 195 191
rect 199 187 205 191
rect -2 183 6 187
rect -2 179 0 183
rect 4 179 8 183
rect 23 179 51 183
rect 55 179 83 183
rect 87 179 99 183
rect 103 179 115 183
rect 119 179 131 183
rect 135 179 163 183
rect 167 179 195 183
rect 199 179 205 183
rect -2 175 6 179
rect -2 171 0 175
rect 4 171 8 175
rect 23 171 51 175
rect 55 171 67 175
rect 71 171 83 175
rect 87 171 99 175
rect 103 171 115 175
rect 119 171 131 175
rect 135 171 163 175
rect 167 171 195 175
rect 199 171 205 175
rect -2 167 6 171
rect -2 163 0 167
rect 4 163 6 167
rect 17 163 35 167
rect 39 163 43 167
rect 47 163 51 167
rect 55 163 59 167
rect 63 163 67 167
rect 71 163 75 167
rect 79 163 83 167
rect 87 163 91 167
rect 95 163 99 167
rect 103 163 107 167
rect 111 163 115 167
rect 119 163 123 167
rect 127 163 131 167
rect 135 163 139 167
rect 143 163 147 167
rect 151 163 155 167
rect 159 163 163 167
rect 167 163 171 167
rect 175 163 179 167
rect 183 163 187 167
rect 191 163 195 167
rect 199 163 205 167
rect -2 159 6 163
rect -2 155 0 159
rect 4 155 8 159
rect 23 155 35 159
rect 39 155 51 159
rect 55 155 67 159
rect 71 155 83 159
rect 87 155 115 159
rect 119 155 131 159
rect 135 155 163 159
rect 167 155 179 159
rect 183 155 205 159
rect -2 151 6 155
rect -2 147 0 151
rect 4 147 8 151
rect 23 147 35 151
rect 39 147 51 151
rect 55 147 67 151
rect 71 147 99 151
rect 103 147 115 151
rect 119 147 131 151
rect 135 147 163 151
rect 167 147 179 151
rect 183 147 205 151
rect -2 143 6 147
rect -2 139 0 143
rect 4 139 6 143
rect 17 139 35 143
rect 39 139 43 143
rect 47 139 51 143
rect 55 139 59 143
rect 63 139 67 143
rect 71 139 75 143
rect 79 139 83 143
rect 87 139 91 143
rect 95 139 99 143
rect 103 139 107 143
rect 111 139 115 143
rect 119 139 123 143
rect 127 139 131 143
rect 135 139 139 143
rect 143 139 147 143
rect 151 139 155 143
rect 159 139 163 143
rect 167 139 171 143
rect 175 139 179 143
rect 183 139 187 143
rect 191 139 195 143
rect 199 139 205 143
rect -2 135 6 139
rect -2 131 0 135
rect 4 131 8 135
rect 23 131 35 135
rect 39 131 51 135
rect 55 131 67 135
rect 71 131 83 135
rect 87 131 99 135
rect 103 131 115 135
rect 119 131 131 135
rect 135 131 163 135
rect 167 131 179 135
rect 183 131 205 135
rect -2 127 6 131
rect -2 123 0 127
rect 4 123 8 127
rect 23 123 51 127
rect 55 123 83 127
rect 87 123 99 127
rect 103 123 115 127
rect 119 123 131 127
rect 135 123 163 127
rect 167 123 179 127
rect 183 123 205 127
rect -2 119 6 123
rect -2 115 0 119
rect 4 115 6 119
rect 17 115 35 119
rect 39 115 43 119
rect 47 115 51 119
rect 55 115 59 119
rect 63 115 67 119
rect 71 115 75 119
rect 79 115 83 119
rect 87 115 91 119
rect 95 115 99 119
rect 103 115 107 119
rect 111 115 115 119
rect 119 115 123 119
rect 127 115 131 119
rect 135 115 139 119
rect 143 115 147 119
rect 151 115 155 119
rect 159 115 163 119
rect 167 115 171 119
rect 175 115 179 119
rect 183 115 187 119
rect 191 115 195 119
rect 199 115 205 119
rect -2 111 6 115
rect -2 107 0 111
rect 4 107 8 111
rect 23 107 51 111
rect 55 107 67 111
rect 71 107 83 111
rect 87 107 99 111
rect 103 107 115 111
rect 119 107 131 111
rect 135 107 163 111
rect 167 107 179 111
rect 183 107 205 111
rect -2 103 6 107
rect -2 99 0 103
rect 4 99 8 103
rect 23 99 131 103
rect 135 99 147 103
rect 151 99 179 103
rect 183 99 195 103
rect 199 99 205 103
rect -2 95 6 99
rect -2 91 0 95
rect 4 91 6 95
rect 17 91 35 95
rect 39 91 43 95
rect 47 91 51 95
rect 55 91 59 95
rect 63 91 67 95
rect 71 91 75 95
rect 79 91 83 95
rect 87 91 91 95
rect 95 91 99 95
rect 103 91 107 95
rect 111 91 115 95
rect 119 91 123 95
rect 127 91 131 95
rect 135 91 139 95
rect 143 91 147 95
rect 151 91 155 95
rect 159 91 163 95
rect 167 91 171 95
rect 175 91 179 95
rect 183 91 187 95
rect 191 91 195 95
rect 199 91 205 95
rect -2 87 6 91
rect -2 83 0 87
rect 4 83 8 87
rect 23 83 131 87
rect 135 83 147 87
rect 151 83 179 87
rect 183 83 205 87
rect -2 79 6 83
rect -2 75 0 79
rect 4 75 8 79
rect 23 75 131 79
rect 135 75 147 79
rect 151 75 163 79
rect 167 75 195 79
rect 199 75 205 79
rect -2 71 6 75
rect -2 67 0 71
rect 4 67 6 71
rect 17 67 35 71
rect 39 67 43 71
rect 47 67 51 71
rect 55 67 59 71
rect 63 67 67 71
rect 71 67 75 71
rect 79 67 83 71
rect 87 67 91 71
rect 95 67 99 71
rect 103 67 107 71
rect 111 67 115 71
rect 119 67 123 71
rect 127 67 131 71
rect 135 67 139 71
rect 143 67 147 71
rect 151 67 155 71
rect 159 67 163 71
rect 167 67 171 71
rect 175 67 179 71
rect 183 67 187 71
rect 191 67 195 71
rect 199 67 205 71
rect -2 63 6 67
rect -2 59 0 63
rect 4 59 8 63
rect 23 59 131 63
rect 135 59 147 63
rect 151 59 163 63
rect 167 59 179 63
rect 183 59 205 63
rect -2 4 6 59
rect 33 53 211 55
rect 33 49 35 53
rect 39 49 51 53
rect 55 49 67 53
rect 71 49 83 53
rect 87 49 99 53
rect 103 49 115 53
rect 119 49 131 53
rect 135 49 147 53
rect 151 49 163 53
rect 167 49 179 53
rect 183 49 205 53
rect 209 49 211 53
rect 215 53 219 231
rect 223 287 227 308
rect 223 263 227 283
rect 223 251 227 259
rect 223 239 227 247
rect 223 227 227 235
rect 223 215 227 223
rect 223 191 227 211
rect 223 167 227 187
rect 223 143 227 163
rect 223 119 227 139
rect 223 95 227 115
rect 223 71 227 91
rect 215 49 216 53
rect 33 47 211 49
rect 35 42 39 47
rect 43 42 47 43
rect 51 42 55 47
rect 59 42 63 43
rect 67 42 71 47
rect 75 42 79 43
rect 83 42 87 47
rect 91 42 95 43
rect 99 42 103 47
rect 107 42 111 43
rect 115 42 119 47
rect 123 42 127 43
rect 131 42 135 47
rect 139 42 143 43
rect 147 42 151 47
rect 155 42 159 43
rect 163 42 167 47
rect 171 42 175 43
rect 179 42 183 47
rect 187 42 191 43
rect 43 34 47 38
rect 59 34 63 38
rect 75 34 79 38
rect 91 34 95 38
rect 107 34 111 38
rect 123 34 127 38
rect 139 34 143 38
rect 155 34 159 38
rect 171 34 175 38
rect 187 34 191 38
rect 215 42 219 43
rect 223 42 227 67
rect 231 259 235 303
rect 231 53 235 255
rect 234 49 235 53
rect 239 259 243 303
rect 239 53 243 255
rect 247 287 251 308
rect 247 275 251 283
rect 247 263 251 271
rect 247 251 251 259
rect 247 239 251 247
rect 247 215 251 235
rect 247 191 251 211
rect 247 167 251 187
rect 247 143 251 163
rect 247 119 251 139
rect 247 107 251 115
rect 247 95 251 103
rect 247 83 251 91
rect 247 71 251 79
rect 247 59 251 67
rect 239 49 240 53
rect 231 42 235 43
rect 43 30 46 34
rect 59 30 62 34
rect 75 30 78 34
rect 91 30 94 34
rect 107 30 110 34
rect 123 30 126 34
rect 139 30 142 34
rect 155 30 158 34
rect 171 30 174 34
rect 187 30 190 34
rect 35 17 39 18
rect 43 17 47 30
rect 51 17 55 18
rect 59 17 63 30
rect 67 17 71 18
rect 75 17 79 30
rect 83 17 87 18
rect 91 17 95 30
rect 99 17 103 18
rect 107 17 111 30
rect 115 17 119 18
rect 123 17 127 30
rect 131 17 135 18
rect 139 17 143 30
rect 147 17 151 18
rect 155 17 159 30
rect 163 17 167 18
rect 171 17 175 30
rect 179 17 183 18
rect 187 17 191 30
rect 215 26 219 38
rect 215 17 219 22
rect 231 26 235 38
rect 223 17 227 18
rect 231 17 235 22
rect 239 42 243 43
rect 247 42 251 55
rect 255 267 259 303
rect 255 99 259 263
rect 255 91 259 95
rect 255 75 259 87
rect 255 67 259 71
rect 255 53 259 63
rect 258 49 259 53
rect 263 99 267 303
rect 263 53 267 95
rect 271 287 275 308
rect 271 263 275 283
rect 271 239 275 259
rect 271 215 275 235
rect 271 191 275 211
rect 271 167 275 187
rect 271 143 275 163
rect 271 119 275 139
rect 271 107 275 115
rect 271 95 275 103
rect 271 83 275 91
rect 271 71 275 79
rect 263 49 264 53
rect 255 42 259 43
rect 239 26 243 38
rect 239 17 243 22
rect 255 26 259 38
rect 247 17 251 18
rect 255 17 259 22
rect 263 42 267 43
rect 271 42 275 67
rect 279 91 283 303
rect 279 53 283 87
rect 282 49 283 53
rect 287 75 291 303
rect 287 53 291 71
rect 295 287 299 308
rect 295 263 299 283
rect 295 239 299 259
rect 295 215 299 235
rect 295 191 299 211
rect 295 167 299 187
rect 295 143 299 163
rect 295 119 299 139
rect 295 95 299 115
rect 295 83 299 91
rect 295 71 299 79
rect 295 59 299 67
rect 287 49 288 53
rect 279 42 283 43
rect 263 26 267 38
rect 263 17 267 22
rect 279 26 283 38
rect 271 17 275 18
rect 279 17 283 22
rect 287 42 291 43
rect 295 42 299 55
rect 303 67 307 303
rect 303 53 307 63
rect 306 49 307 53
rect 311 187 315 303
rect 311 171 315 183
rect 311 163 315 167
rect 311 147 315 159
rect 311 139 315 143
rect 311 123 315 135
rect 311 115 315 119
rect 311 53 315 111
rect 319 287 323 308
rect 319 263 323 283
rect 319 239 323 259
rect 319 215 323 235
rect 319 191 323 211
rect 319 179 323 187
rect 319 167 323 175
rect 319 155 323 163
rect 319 143 323 151
rect 319 131 323 139
rect 319 119 323 127
rect 319 107 323 115
rect 319 95 323 103
rect 319 83 323 91
rect 319 71 323 79
rect 319 59 323 67
rect 311 49 312 53
rect 303 42 307 43
rect 287 26 291 38
rect 287 17 291 22
rect 303 26 307 38
rect 295 17 299 18
rect 303 17 307 22
rect 311 42 315 43
rect 319 42 323 55
rect 327 163 331 303
rect 327 147 331 159
rect 327 139 331 143
rect 327 123 331 135
rect 327 115 331 119
rect 327 99 331 111
rect 327 91 331 95
rect 327 75 331 87
rect 327 67 331 71
rect 327 53 331 63
rect 330 49 331 53
rect 335 267 339 303
rect 335 53 339 263
rect 343 287 347 308
rect 343 275 347 283
rect 343 263 347 271
rect 343 251 347 259
rect 343 239 347 247
rect 343 215 347 235
rect 343 191 347 211
rect 343 167 347 187
rect 343 143 347 163
rect 343 119 347 139
rect 343 95 347 115
rect 343 71 347 91
rect 335 49 336 53
rect 327 42 331 43
rect 311 26 315 38
rect 311 17 315 22
rect 327 26 331 38
rect 319 17 323 18
rect 327 17 331 22
rect 335 42 339 43
rect 343 42 347 67
rect 351 259 355 303
rect 351 53 355 255
rect 354 49 355 53
rect 359 243 363 303
rect 359 53 363 239
rect 367 287 371 308
rect 367 275 371 283
rect 367 263 371 271
rect 367 251 371 259
rect 367 239 371 247
rect 367 215 371 235
rect 367 203 371 211
rect 367 191 371 199
rect 367 167 371 187
rect 367 143 371 163
rect 367 119 371 139
rect 367 95 371 115
rect 367 71 371 91
rect 359 49 360 53
rect 351 42 355 43
rect 335 26 339 38
rect 335 17 339 22
rect 351 26 355 38
rect 343 17 347 18
rect 351 17 355 22
rect 359 42 363 43
rect 367 42 371 67
rect 375 283 379 303
rect 375 243 379 279
rect 375 211 379 239
rect 375 53 379 207
rect 378 49 379 53
rect 383 219 387 303
rect 383 195 387 215
rect 383 53 387 191
rect 391 287 395 308
rect 391 263 395 283
rect 391 239 395 259
rect 391 227 395 235
rect 391 215 395 223
rect 391 203 395 211
rect 391 191 395 199
rect 391 167 395 187
rect 391 143 395 163
rect 391 119 395 139
rect 391 95 395 115
rect 391 71 395 91
rect 383 49 384 53
rect 375 42 379 43
rect 359 26 363 38
rect 359 17 363 22
rect 375 26 379 38
rect 367 17 371 18
rect 375 17 379 22
rect 383 42 387 43
rect 391 42 395 67
rect 399 211 403 303
rect 399 53 403 207
rect 402 49 403 53
rect 407 259 411 303
rect 407 235 411 255
rect 407 187 411 231
rect 407 171 411 183
rect 407 53 411 167
rect 415 287 419 308
rect 415 263 419 283
rect 415 251 419 259
rect 415 239 419 247
rect 415 227 419 235
rect 415 215 419 223
rect 415 191 419 211
rect 415 179 419 187
rect 415 167 419 175
rect 415 143 419 163
rect 415 119 419 139
rect 415 95 419 115
rect 415 71 419 91
rect 407 49 408 53
rect 399 42 403 43
rect 383 26 387 38
rect 383 17 387 22
rect 399 26 403 38
rect 391 17 395 18
rect 399 17 403 22
rect 407 42 411 43
rect 415 42 419 67
rect 423 219 427 303
rect 423 53 427 215
rect 426 49 427 53
rect 431 195 435 303
rect 431 99 435 191
rect 431 91 435 95
rect 431 75 435 87
rect 431 67 435 71
rect 431 53 435 63
rect 439 287 443 308
rect 439 263 443 283
rect 439 239 443 259
rect 439 227 443 235
rect 439 215 443 223
rect 439 203 443 211
rect 439 191 443 199
rect 439 179 443 187
rect 439 167 443 175
rect 439 155 443 163
rect 439 143 443 151
rect 439 131 443 139
rect 439 119 443 127
rect 439 107 443 115
rect 439 95 443 103
rect 439 83 443 91
rect 439 71 443 79
rect 439 59 443 67
rect 431 49 432 53
rect 423 42 427 43
rect 407 26 411 38
rect 407 17 411 22
rect 423 26 427 38
rect 415 17 419 18
rect 423 17 427 22
rect 431 42 435 43
rect 439 42 443 55
rect 447 235 451 303
rect 447 187 451 231
rect 447 163 451 183
rect 447 147 451 159
rect 447 139 451 143
rect 447 53 451 135
rect 450 49 451 53
rect 455 195 459 303
rect 455 171 459 191
rect 455 163 459 167
rect 455 123 459 159
rect 455 115 459 119
rect 455 99 459 111
rect 455 53 459 95
rect 463 287 467 308
rect 463 263 467 283
rect 463 239 467 259
rect 463 227 467 235
rect 463 215 467 223
rect 463 203 467 211
rect 463 191 467 199
rect 463 179 467 187
rect 463 167 467 175
rect 463 155 467 163
rect 463 143 467 151
rect 463 131 467 139
rect 463 119 467 127
rect 463 107 467 115
rect 463 95 467 103
rect 463 83 467 91
rect 463 71 467 79
rect 455 49 456 53
rect 447 42 451 43
rect 431 26 435 38
rect 431 17 435 22
rect 447 26 451 38
rect 439 17 443 18
rect 447 17 451 22
rect 455 42 459 43
rect 463 42 467 67
rect 471 235 475 303
rect 471 195 475 231
rect 471 171 475 191
rect 471 147 475 167
rect 471 91 475 143
rect 471 75 475 87
rect 471 53 475 71
rect 474 49 475 53
rect 479 195 483 303
rect 479 147 483 191
rect 479 139 483 143
rect 479 123 483 135
rect 479 115 483 119
rect 479 91 483 111
rect 479 67 483 87
rect 479 53 483 63
rect 487 287 491 308
rect 487 263 491 283
rect 487 239 491 259
rect 487 215 491 235
rect 487 203 491 211
rect 487 191 491 199
rect 487 167 491 187
rect 487 155 491 163
rect 487 143 491 151
rect 487 131 491 139
rect 487 119 491 127
rect 487 107 491 115
rect 487 95 491 103
rect 487 83 491 91
rect 487 71 491 79
rect 487 59 491 67
rect 479 49 480 53
rect 471 42 475 43
rect 455 26 459 38
rect 455 17 459 22
rect 471 26 475 38
rect 463 17 467 18
rect 471 17 475 22
rect 479 42 483 43
rect 487 42 491 55
rect 479 26 483 38
rect 479 17 483 22
rect 487 17 491 18
rect 35 4 39 8
rect 51 4 55 8
rect 67 4 71 8
rect 83 4 87 8
rect 99 4 103 8
rect 115 4 119 8
rect 131 4 135 8
rect 147 4 151 8
rect 163 4 167 8
rect 179 4 183 8
rect 223 4 227 8
rect 247 4 251 8
rect 271 4 275 8
rect 295 4 299 8
rect 319 4 323 8
rect 343 4 347 8
rect 367 4 371 8
rect 391 4 395 8
rect 415 4 419 8
rect 439 4 443 8
rect 463 4 467 8
rect 487 4 491 8
rect -2 2 493 4
rect -2 -2 0 2
rect 4 -2 35 2
rect 39 -2 43 2
rect 47 -2 51 2
rect 55 -2 59 2
rect 63 -2 67 2
rect 71 -2 75 2
rect 79 -2 83 2
rect 87 -2 91 2
rect 95 -2 99 2
rect 103 -2 107 2
rect 111 -2 115 2
rect 119 -2 123 2
rect 127 -2 131 2
rect 135 -2 139 2
rect 143 -2 147 2
rect 151 -2 155 2
rect 159 -2 163 2
rect 167 -2 171 2
rect 175 -2 179 2
rect 183 -2 187 2
rect 191 -2 215 2
rect 219 -2 223 2
rect 227 -2 231 2
rect 235 -2 239 2
rect 243 -2 247 2
rect 251 -2 255 2
rect 259 -2 263 2
rect 267 -2 271 2
rect 275 -2 279 2
rect 283 -2 287 2
rect 291 -2 295 2
rect 299 -2 303 2
rect 307 -2 311 2
rect 315 -2 319 2
rect 323 -2 327 2
rect 331 -2 335 2
rect 339 -2 343 2
rect 347 -2 351 2
rect 355 -2 359 2
rect 363 -2 367 2
rect 371 -2 375 2
rect 379 -2 383 2
rect 387 -2 391 2
rect 395 -2 399 2
rect 403 -2 407 2
rect 411 -2 415 2
rect 419 -2 423 2
rect 427 -2 431 2
rect 435 -2 439 2
rect 443 -2 447 2
rect 451 -2 455 2
rect 459 -2 463 2
rect 467 -2 471 2
rect 475 -2 479 2
rect 483 -2 487 2
rect 491 -2 493 2
rect -2 -4 493 -2
<< m2contact >>
rect 205 334 209 338
rect 223 334 227 338
rect 247 334 251 338
rect 271 334 275 338
rect 295 334 299 338
rect 319 334 323 338
rect 343 334 347 338
rect 367 334 371 338
rect 391 334 395 338
rect 415 334 419 338
rect 439 334 443 338
rect 463 334 467 338
rect 487 334 491 338
rect 223 308 227 312
rect 205 283 209 287
rect 205 259 209 263
rect 205 235 209 239
rect 205 211 209 215
rect 205 187 209 191
rect 205 163 209 167
rect 205 139 209 143
rect 205 115 209 119
rect 205 91 209 95
rect 205 67 209 71
rect 205 49 209 53
rect 247 308 251 312
rect 271 308 275 312
rect 35 22 39 26
rect 51 22 55 26
rect 67 22 71 26
rect 83 22 84 26
rect 84 22 87 26
rect 99 22 100 26
rect 100 22 103 26
rect 115 22 116 26
rect 116 22 119 26
rect 131 22 132 26
rect 132 22 135 26
rect 147 22 148 26
rect 148 22 151 26
rect 163 22 164 26
rect 164 22 167 26
rect 179 22 180 26
rect 180 22 183 26
rect 215 22 219 26
rect 231 22 235 26
rect 295 308 299 312
rect 239 22 243 26
rect 255 22 259 26
rect 319 308 323 312
rect 263 22 267 26
rect 279 22 283 26
rect 343 308 347 312
rect 287 22 291 26
rect 303 22 307 26
rect 367 308 371 312
rect 311 22 315 26
rect 327 22 331 26
rect 391 308 395 312
rect 335 22 339 26
rect 351 22 355 26
rect 415 308 419 312
rect 359 22 363 26
rect 375 22 379 26
rect 439 308 443 312
rect 383 22 387 26
rect 399 22 403 26
rect 463 308 467 312
rect 407 22 411 26
rect 423 22 427 26
rect 487 308 491 312
rect 431 22 435 26
rect 447 22 451 26
rect 455 22 459 26
rect 471 22 475 26
rect 479 22 483 26
rect 0 -2 4 2
<< metal2 >>
rect 203 338 211 340
rect 203 334 205 338
rect 209 334 211 338
rect 203 287 211 334
rect 223 312 227 334
rect 247 312 251 334
rect 271 312 275 334
rect 295 312 299 334
rect 319 312 323 334
rect 343 312 347 334
rect 367 312 371 334
rect 391 312 395 334
rect 415 312 419 334
rect 439 312 443 334
rect 463 312 467 334
rect 487 312 491 334
rect 203 283 205 287
rect 209 283 211 287
rect 203 263 211 283
rect 203 259 205 263
rect 209 259 211 263
rect 203 239 211 259
rect 203 235 205 239
rect 209 235 211 239
rect 203 215 211 235
rect 203 211 205 215
rect 209 211 211 215
rect 203 191 211 211
rect 203 187 205 191
rect 209 187 211 191
rect 203 167 211 187
rect 203 163 205 167
rect 209 163 211 167
rect 203 143 211 163
rect 203 139 205 143
rect 209 139 211 143
rect 203 119 211 139
rect 203 115 205 119
rect 209 115 211 119
rect 203 95 211 115
rect 203 91 205 95
rect 209 91 211 95
rect 203 71 211 91
rect 203 67 205 71
rect 209 67 211 71
rect 203 53 211 67
rect 203 49 205 53
rect 209 49 211 53
rect 203 47 211 49
<< labels >>
rlabel m2contact 37 24 37 24 1 in_9_
rlabel m2contact 69 24 69 24 1 in_7_
rlabel m2contact 53 24 53 24 1 in_8_
rlabel m2contact 85 24 85 24 1 in_6_
rlabel m2contact 101 24 101 24 1 in_5_
rlabel m2contact 117 24 117 24 1 in_4_
rlabel m2contact 133 24 133 24 1 in_3_
rlabel m2contact 149 24 149 24 1 in_2_
rlabel m2contact 165 24 165 24 1 in_1_
rlabel metal1 105 324 105 324 1 Vdd!
rlabel metal1 219 336 219 336 5 Gnd!
rlabel metal1 481 28 481 28 1 out_0_
rlabel metal1 473 28 473 28 1 out_1_
rlabel metal1 457 28 457 28 1 out_2_
rlabel metal1 449 28 449 28 1 out_3_
rlabel metal1 433 28 433 28 1 out_4_
rlabel metal1 425 28 425 28 1 out_5_
rlabel metal1 409 28 409 28 1 out_6_
rlabel metal1 401 28 401 28 1 out_7_
rlabel metal1 385 28 385 28 1 out_8_
rlabel metal1 377 28 377 28 1 out_9_
rlabel metal1 361 28 361 28 1 out_10_
rlabel metal1 353 28 353 28 1 out_11_
rlabel metal1 329 28 329 28 1 out_13_
rlabel metal1 337 28 337 28 1 out_12_
rlabel metal1 313 28 313 28 1 out_14_
rlabel metal1 305 28 305 28 1 out_15_
rlabel metal1 289 28 289 28 1 out_16_
rlabel metal1 281 28 281 28 1 out_17_
rlabel metal1 265 28 265 28 1 out_18_
rlabel metal1 257 28 257 28 1 out_18_
rlabel metal1 257 28 257 28 1 out_19_
rlabel metal1 241 28 241 28 1 out_20_
rlabel metal1 233 28 233 28 1 out_21_
rlabel metal1 217 29 217 29 1 out_22_
<< end >>
