magic
tech scmos
timestamp 1271709725
<< nwell >>
rect 20 740 280 1000
rect 17 429 283 653
rect -3 248 303 330
rect -3 11 11 248
rect 289 11 303 248
rect -3 -3 303 11
<< pwell >>
rect -3 656 303 673
rect -3 426 14 656
rect 286 426 303 656
rect -3 340 303 426
rect 11 11 289 248
<< ntransistor >>
rect 38 216 138 219
rect 162 216 262 219
rect 38 171 138 174
rect 38 150 138 153
rect 162 171 262 174
rect 162 150 262 153
rect 38 106 138 109
rect 38 85 138 88
rect 162 106 262 109
rect 162 85 262 88
rect 38 41 138 44
rect 162 41 262 44
<< ptransistor >>
rect 38 626 138 629
rect 162 626 262 629
rect 38 582 138 585
rect 38 562 138 565
rect 162 582 262 585
rect 162 562 262 565
rect 38 518 138 521
rect 38 497 138 500
rect 162 518 262 521
rect 162 497 262 500
rect 38 453 138 456
rect 162 453 262 456
<< ndiffusion >>
rect 38 227 138 228
rect 38 223 41 227
rect 95 223 138 227
rect 38 219 138 223
rect 162 227 262 228
rect 162 223 205 227
rect 259 223 262 227
rect 162 219 262 223
rect 38 200 138 216
rect 38 196 56 200
rect 120 196 138 200
rect 38 194 138 196
rect 38 190 56 194
rect 120 190 138 194
rect 38 174 138 190
rect 38 167 138 171
rect 38 163 41 167
rect 120 163 138 167
rect 38 161 138 163
rect 38 157 41 161
rect 120 157 138 161
rect 38 153 138 157
rect 38 134 138 150
rect 38 125 56 134
rect 120 125 138 134
rect 38 109 138 125
rect 162 200 262 216
rect 162 196 180 200
rect 244 196 262 200
rect 162 194 262 196
rect 162 190 180 194
rect 244 190 262 194
rect 162 174 262 190
rect 162 167 262 171
rect 162 163 180 167
rect 259 163 262 167
rect 162 161 262 163
rect 162 157 180 161
rect 259 157 262 161
rect 162 153 262 157
rect 38 102 138 106
rect 38 98 41 102
rect 120 98 138 102
rect 38 96 138 98
rect 38 92 41 96
rect 120 92 138 96
rect 38 88 138 92
rect 38 69 138 85
rect 38 60 56 69
rect 120 60 138 69
rect 38 44 138 60
rect 162 134 262 150
rect 162 125 180 134
rect 244 125 262 134
rect 162 109 262 125
rect 162 102 262 106
rect 162 98 180 102
rect 259 98 262 102
rect 162 96 262 98
rect 162 92 180 96
rect 259 92 262 96
rect 162 88 262 92
rect 162 69 262 85
rect 162 60 180 69
rect 244 60 262 69
rect 162 44 262 60
rect 38 37 138 41
rect 38 33 41 37
rect 95 33 138 37
rect 38 32 138 33
rect 162 37 262 41
rect 162 33 205 37
rect 259 33 262 37
rect 162 32 262 33
<< pdiffusion >>
rect 38 636 138 638
rect 38 632 41 636
rect 120 632 138 636
rect 38 629 138 632
rect 38 610 138 626
rect 38 601 56 610
rect 120 601 138 610
rect 38 585 138 601
rect 162 636 262 638
rect 162 632 180 636
rect 259 632 262 636
rect 162 629 262 632
rect 38 578 138 582
rect 38 569 41 578
rect 120 569 138 578
rect 38 565 138 569
rect 38 546 138 562
rect 38 537 56 546
rect 120 537 138 546
rect 38 521 138 537
rect 162 610 262 626
rect 162 601 180 610
rect 244 601 262 610
rect 162 585 262 601
rect 162 578 262 582
rect 162 569 180 578
rect 259 569 262 578
rect 162 565 262 569
rect 38 514 138 518
rect 38 510 41 514
rect 120 510 138 514
rect 38 508 138 510
rect 38 504 41 508
rect 120 504 138 508
rect 38 500 138 504
rect 38 481 138 497
rect 38 472 56 481
rect 120 472 138 481
rect 38 456 138 472
rect 162 546 262 562
rect 162 537 180 546
rect 244 537 262 546
rect 162 521 262 537
rect 162 514 262 518
rect 162 510 180 514
rect 259 510 262 514
rect 162 508 262 510
rect 162 504 180 508
rect 259 504 262 508
rect 162 500 262 504
rect 38 449 138 453
rect 38 445 41 449
rect 120 445 138 449
rect 38 444 138 445
rect 162 481 262 497
rect 162 472 180 481
rect 244 472 262 481
rect 162 456 262 472
rect 162 449 262 453
rect 162 445 180 449
rect 259 445 262 449
rect 162 444 262 445
<< ndcontact >>
rect 41 223 95 227
rect 205 223 259 227
rect 56 196 120 200
rect 56 190 120 194
rect 41 163 120 167
rect 41 157 120 161
rect 56 125 120 134
rect 180 196 244 200
rect 180 190 244 194
rect 180 163 259 167
rect 180 157 259 161
rect 41 98 120 102
rect 41 92 120 96
rect 56 60 120 69
rect 180 125 244 134
rect 180 98 259 102
rect 180 92 259 96
rect 180 60 244 69
rect 41 33 95 37
rect 205 33 259 37
<< pdcontact >>
rect 41 632 120 636
rect 56 601 120 610
rect 180 632 259 636
rect 41 569 120 578
rect 56 537 120 546
rect 180 601 244 610
rect 180 569 259 578
rect 41 510 120 514
rect 41 504 120 508
rect 56 472 120 481
rect 180 537 244 546
rect 180 510 259 514
rect 180 504 259 508
rect 41 445 120 449
rect 180 472 244 481
rect 180 445 259 449
<< psubstratepdiff >>
rect 0 669 300 670
rect 0 660 1 669
rect 99 660 201 669
rect 299 660 300 669
rect 0 659 300 660
rect 0 658 11 659
rect 0 424 1 658
rect 10 424 11 658
rect 289 658 300 659
rect 0 423 11 424
rect 289 424 290 658
rect 299 424 300 658
rect 289 423 300 424
rect 0 418 300 423
rect 0 414 3 418
rect 96 414 143 418
rect 157 414 204 418
rect 298 414 300 418
rect 0 408 300 414
rect 0 404 3 408
rect 96 404 143 408
rect 157 404 204 408
rect 298 404 300 408
rect 0 398 300 404
rect 0 394 3 398
rect 96 394 143 398
rect 157 394 204 398
rect 298 394 300 398
rect 0 388 300 394
rect 0 384 3 388
rect 96 384 143 388
rect 157 384 204 388
rect 298 384 300 388
rect 0 378 300 384
rect 0 374 3 378
rect 96 374 143 378
rect 157 374 204 378
rect 298 374 300 378
rect 0 368 300 374
rect 0 364 3 368
rect 96 364 143 368
rect 157 364 204 368
rect 298 364 300 368
rect 0 358 300 364
rect 0 354 3 358
rect 96 354 143 358
rect 157 354 204 358
rect 298 354 300 358
rect 0 348 300 354
rect 0 344 3 348
rect 96 344 143 348
rect 157 344 204 348
rect 298 344 300 348
rect 0 343 300 344
rect 14 244 286 245
rect 14 241 202 244
rect 14 237 19 241
rect 98 237 202 241
rect 14 235 202 237
rect 281 235 286 244
rect 14 233 286 235
rect 14 29 24 233
rect 28 230 39 233
rect 28 30 30 230
rect 38 229 39 230
rect 98 230 202 233
rect 98 229 138 230
rect 38 228 138 229
rect 142 223 158 230
rect 142 219 145 223
rect 154 219 158 223
rect 162 229 202 230
rect 261 230 277 233
rect 261 229 262 230
rect 162 228 262 229
rect 142 215 158 219
rect 142 211 145 215
rect 154 211 158 215
rect 142 207 158 211
rect 142 203 145 207
rect 154 203 158 207
rect 142 135 158 203
rect 142 131 145 135
rect 154 131 158 135
rect 142 127 158 131
rect 142 123 145 127
rect 154 123 158 127
rect 142 63 158 123
rect 142 59 145 63
rect 154 59 158 63
rect 142 55 158 59
rect 142 51 145 55
rect 154 51 158 55
rect 142 47 158 51
rect 142 43 145 47
rect 154 43 158 47
rect 38 30 138 32
rect 142 39 158 43
rect 142 35 145 39
rect 154 35 158 39
rect 142 30 158 35
rect 162 30 262 32
rect 270 30 277 230
rect 28 29 277 30
rect 281 29 286 233
rect 14 27 286 29
rect 14 23 19 27
rect 98 23 202 27
rect 281 23 286 27
rect 14 14 286 23
<< nsubstratendiff >>
rect 20 649 280 650
rect 20 445 26 649
rect 30 647 270 649
rect 30 643 36 647
rect 120 643 180 647
rect 264 643 270 647
rect 30 640 270 643
rect 36 638 138 640
rect 142 615 158 640
rect 162 638 264 640
rect 142 611 143 615
rect 157 611 158 615
rect 142 605 158 611
rect 142 601 143 605
rect 157 601 158 605
rect 142 595 158 601
rect 142 591 143 595
rect 157 591 158 595
rect 142 551 158 591
rect 142 547 143 551
rect 157 547 158 551
rect 142 541 158 547
rect 142 537 143 541
rect 157 537 158 541
rect 142 531 158 537
rect 142 527 143 531
rect 157 527 158 531
rect 142 486 158 527
rect 142 482 143 486
rect 157 482 158 486
rect 142 476 158 482
rect 142 472 143 476
rect 157 472 158 476
rect 142 466 158 472
rect 142 462 143 466
rect 157 462 158 466
rect 20 442 30 445
rect 38 442 138 444
rect 142 442 158 462
rect 162 442 262 444
rect 274 445 280 649
rect 270 442 280 445
rect 20 441 280 442
rect 20 432 21 441
rect 120 432 180 441
rect 279 432 280 441
rect 0 326 300 327
rect 0 322 2 326
rect 96 322 143 326
rect 157 322 204 326
rect 298 322 300 326
rect 0 316 300 322
rect 0 312 2 316
rect 96 312 143 316
rect 157 312 204 316
rect 298 312 300 316
rect 0 306 300 312
rect 0 302 2 306
rect 96 302 143 306
rect 157 302 204 306
rect 298 302 300 306
rect 0 296 300 302
rect 0 292 2 296
rect 96 292 143 296
rect 157 292 204 296
rect 298 292 300 296
rect 0 286 300 292
rect 0 282 2 286
rect 96 282 143 286
rect 157 282 204 286
rect 298 282 300 286
rect 0 276 300 282
rect 0 272 2 276
rect 96 272 143 276
rect 157 272 204 276
rect 298 272 300 276
rect 0 266 300 272
rect 0 262 2 266
rect 96 262 143 266
rect 157 262 204 266
rect 298 262 300 266
rect 0 256 300 262
rect 0 3 2 256
rect 6 8 8 256
rect 97 252 143 256
rect 157 252 203 256
rect 292 8 294 256
rect 6 7 294 8
rect 6 3 8 7
rect 92 3 203 7
rect 292 3 294 7
rect 298 3 300 256
rect 0 0 300 3
<< psubstratepcontact >>
rect 1 660 99 669
rect 201 660 299 669
rect 1 424 10 658
rect 290 424 299 658
rect 3 414 96 418
rect 143 414 157 418
rect 204 414 298 418
rect 3 404 96 408
rect 143 404 157 408
rect 204 404 298 408
rect 3 394 96 398
rect 143 394 157 398
rect 204 394 298 398
rect 3 384 96 388
rect 143 384 157 388
rect 204 384 298 388
rect 3 374 96 378
rect 143 374 157 378
rect 204 374 298 378
rect 3 364 96 368
rect 143 364 157 368
rect 204 364 298 368
rect 3 354 96 358
rect 143 354 157 358
rect 204 354 298 358
rect 3 344 96 348
rect 143 344 157 348
rect 204 344 298 348
rect 19 237 98 241
rect 202 235 281 244
rect 24 29 28 233
rect 39 229 98 233
rect 145 219 154 223
rect 202 229 261 233
rect 145 211 154 215
rect 145 203 154 207
rect 145 131 154 135
rect 145 123 154 127
rect 145 59 154 63
rect 145 51 154 55
rect 145 43 154 47
rect 145 35 154 39
rect 277 29 281 233
rect 19 23 98 27
rect 202 23 281 27
<< nsubstratencontact >>
rect 26 445 30 649
rect 36 643 120 647
rect 180 643 264 647
rect 143 611 157 615
rect 143 601 157 605
rect 143 591 157 595
rect 143 547 157 551
rect 143 537 157 541
rect 143 527 157 531
rect 143 482 157 486
rect 143 472 157 476
rect 143 462 157 466
rect 270 445 274 649
rect 21 432 120 441
rect 180 432 279 441
rect 2 322 96 326
rect 143 322 157 326
rect 204 322 298 326
rect 2 312 96 316
rect 143 312 157 316
rect 204 312 298 316
rect 2 302 96 306
rect 143 302 157 306
rect 204 302 298 306
rect 2 292 96 296
rect 143 292 157 296
rect 204 292 298 296
rect 2 282 96 286
rect 143 282 157 286
rect 204 282 298 286
rect 2 272 96 276
rect 143 272 157 276
rect 204 272 298 276
rect 2 262 96 266
rect 143 262 157 266
rect 204 262 298 266
rect 2 3 6 256
rect 8 252 97 256
rect 143 252 157 256
rect 203 252 292 256
rect 8 3 92 7
rect 203 3 292 7
rect 294 3 298 256
<< polysilicon >>
rect 31 626 38 629
rect 138 626 140 629
rect 31 457 32 626
rect 36 585 37 626
rect 160 626 162 629
rect 262 626 269 629
rect 36 582 38 585
rect 138 582 140 585
rect 36 565 37 582
rect 36 562 38 565
rect 138 562 140 565
rect 36 521 37 562
rect 263 585 264 626
rect 160 582 162 585
rect 262 582 264 585
rect 263 565 264 582
rect 160 562 162 565
rect 262 562 264 565
rect 36 518 38 521
rect 138 518 140 521
rect 36 500 37 518
rect 36 497 38 500
rect 138 497 140 500
rect 36 457 37 497
rect 31 456 37 457
rect 263 521 264 562
rect 160 518 162 521
rect 262 518 264 521
rect 263 500 264 518
rect 160 497 162 500
rect 262 497 264 500
rect 31 453 38 456
rect 138 453 140 456
rect 263 457 264 497
rect 268 457 269 626
rect 263 456 269 457
rect 160 453 162 456
rect 262 453 269 456
rect 31 217 38 219
rect 31 43 32 217
rect 36 216 38 217
rect 138 216 140 219
rect 36 174 37 216
rect 160 216 162 219
rect 262 217 269 219
rect 262 216 264 217
rect 36 171 38 174
rect 138 171 140 174
rect 36 153 37 171
rect 36 150 38 153
rect 138 150 140 153
rect 36 109 37 150
rect 263 174 264 216
rect 160 171 162 174
rect 262 171 264 174
rect 263 153 264 171
rect 160 150 162 153
rect 262 150 264 153
rect 36 106 38 109
rect 138 106 140 109
rect 36 88 37 106
rect 36 85 38 88
rect 138 85 140 88
rect 36 44 37 85
rect 263 109 264 150
rect 160 106 162 109
rect 262 106 264 109
rect 263 88 264 106
rect 160 85 162 88
rect 262 85 264 88
rect 36 43 38 44
rect 31 41 38 43
rect 138 41 140 44
rect 263 44 264 85
rect 160 41 162 44
rect 262 43 264 44
rect 268 43 269 217
rect 262 41 269 43
<< polycontact >>
rect 32 457 36 626
rect 264 457 268 626
rect 32 43 36 217
rect 264 43 268 217
<< metal1 >>
rect 20 997 280 1000
rect 20 743 23 997
rect 277 743 280 997
rect 20 740 280 743
rect 62 730 238 740
rect 72 720 228 730
rect 82 710 218 720
rect 92 700 208 710
rect 0 669 99 670
rect 0 660 1 669
rect 0 659 99 660
rect 0 658 11 659
rect 0 424 1 658
rect 10 424 11 658
rect 102 653 198 700
rect 201 669 300 670
rect 299 660 300 669
rect 201 659 300 660
rect 289 658 300 659
rect 36 649 120 650
rect 20 445 21 649
rect 25 445 26 649
rect 30 647 120 649
rect 30 643 36 647
rect 30 642 120 643
rect 30 638 36 642
rect 30 636 120 638
rect 30 632 41 636
rect 30 626 120 632
rect 30 457 32 626
rect 36 625 120 626
rect 36 586 39 625
rect 48 621 52 625
rect 116 621 120 625
rect 48 590 51 621
rect 123 618 177 653
rect 180 649 280 650
rect 180 647 270 649
rect 264 643 270 647
rect 180 642 270 643
rect 264 638 270 642
rect 180 636 270 638
rect 259 632 270 636
rect 180 626 270 632
rect 180 625 264 626
rect 180 621 184 625
rect 248 621 252 625
rect 56 610 140 618
rect 120 601 140 610
rect 56 593 140 601
rect 48 586 52 590
rect 116 586 120 590
rect 36 578 120 586
rect 36 569 41 578
rect 36 561 120 569
rect 36 522 39 561
rect 48 557 52 561
rect 116 557 120 561
rect 123 588 140 593
rect 143 610 157 611
rect 143 605 157 606
rect 143 600 157 601
rect 143 595 157 596
rect 160 610 244 618
rect 160 601 180 610
rect 160 593 244 601
rect 160 588 177 593
rect 249 590 252 621
rect 48 526 51 557
rect 123 554 177 588
rect 180 586 184 590
rect 248 586 252 590
rect 261 586 264 625
rect 180 578 264 586
rect 259 569 264 578
rect 180 561 264 569
rect 180 557 184 561
rect 248 557 252 561
rect 56 546 140 554
rect 120 537 140 546
rect 56 529 140 537
rect 48 522 52 526
rect 116 522 120 526
rect 36 514 120 522
rect 36 510 41 514
rect 36 508 120 510
rect 36 504 41 508
rect 36 496 120 504
rect 36 457 39 496
rect 48 492 52 496
rect 116 492 120 496
rect 123 524 140 529
rect 143 546 157 547
rect 143 541 157 542
rect 143 536 157 537
rect 143 531 157 532
rect 160 546 244 554
rect 160 537 180 546
rect 160 529 244 537
rect 160 524 177 529
rect 249 526 252 557
rect 48 461 51 492
rect 123 489 177 524
rect 180 522 184 526
rect 248 522 252 526
rect 261 522 264 561
rect 180 514 264 522
rect 259 510 264 514
rect 180 508 264 510
rect 259 504 264 508
rect 180 496 264 504
rect 180 492 184 496
rect 248 492 252 496
rect 56 481 140 489
rect 120 472 140 481
rect 56 464 140 472
rect 48 457 52 461
rect 116 457 120 461
rect 30 449 120 457
rect 30 445 41 449
rect 20 441 120 445
rect 20 432 21 441
rect 123 459 140 464
rect 143 481 157 482
rect 143 476 157 477
rect 143 471 157 472
rect 143 466 157 467
rect 160 481 244 489
rect 160 472 180 481
rect 160 464 244 472
rect 160 459 177 464
rect 249 461 252 492
rect 123 429 177 459
rect 180 457 184 461
rect 248 457 252 461
rect 261 457 264 496
rect 268 457 270 626
rect 180 449 270 457
rect 259 445 270 449
rect 274 445 275 649
rect 279 445 280 649
rect 180 441 280 445
rect 279 432 280 441
rect 0 423 11 424
rect 102 424 198 429
rect 0 418 99 423
rect 0 414 3 418
rect 96 414 99 418
rect 0 413 99 414
rect 0 409 3 413
rect 96 409 99 413
rect 0 408 99 409
rect 0 404 3 408
rect 96 404 99 408
rect 0 403 99 404
rect 0 399 3 403
rect 96 399 99 403
rect 0 398 99 399
rect 0 394 3 398
rect 96 394 99 398
rect 0 393 99 394
rect 0 389 3 393
rect 96 389 99 393
rect 0 388 99 389
rect 0 384 3 388
rect 96 384 99 388
rect 0 383 99 384
rect 0 379 3 383
rect 96 379 99 383
rect 0 378 99 379
rect 0 374 3 378
rect 96 374 99 378
rect 0 373 99 374
rect 0 369 3 373
rect 96 369 99 373
rect 0 368 99 369
rect 0 364 3 368
rect 96 364 99 368
rect 0 363 99 364
rect 0 359 3 363
rect 96 359 99 363
rect 0 358 99 359
rect 0 354 3 358
rect 96 354 99 358
rect 0 353 99 354
rect 0 349 3 353
rect 96 349 99 353
rect 0 348 99 349
rect 0 344 3 348
rect 96 344 99 348
rect 102 340 140 424
rect 143 418 157 421
rect 143 413 157 414
rect 143 408 157 409
rect 143 403 157 404
rect 143 398 157 399
rect 143 393 157 394
rect 143 388 157 389
rect 143 383 157 384
rect 143 378 157 379
rect 143 373 157 374
rect 143 368 157 369
rect 143 363 157 364
rect 143 358 157 359
rect 143 353 157 354
rect 143 348 157 349
rect 160 340 198 424
rect 289 424 290 658
rect 299 424 300 658
rect 289 419 300 424
rect 201 418 300 419
rect 201 414 204 418
rect 298 414 300 418
rect 201 413 300 414
rect 201 409 204 413
rect 298 409 300 413
rect 201 408 300 409
rect 201 404 204 408
rect 298 404 300 408
rect 201 403 300 404
rect 201 399 204 403
rect 298 399 300 403
rect 201 398 300 399
rect 201 394 204 398
rect 298 394 300 398
rect 201 393 300 394
rect 201 389 204 393
rect 298 389 300 393
rect 201 388 300 389
rect 201 384 204 388
rect 298 384 300 388
rect 201 383 300 384
rect 201 379 204 383
rect 298 379 300 383
rect 201 378 300 379
rect 201 374 204 378
rect 298 374 300 378
rect 201 373 300 374
rect 201 369 204 373
rect 298 369 300 373
rect 201 368 300 369
rect 201 364 204 368
rect 298 364 300 368
rect 201 363 300 364
rect 201 359 204 363
rect 298 359 300 363
rect 201 358 300 359
rect 201 354 204 358
rect 298 354 300 358
rect 201 353 300 354
rect 201 349 204 353
rect 298 349 300 353
rect 201 348 300 349
rect 201 344 204 348
rect 298 344 300 348
rect 102 329 198 340
rect 0 322 2 326
rect 96 322 99 326
rect 0 321 99 322
rect 0 317 2 321
rect 96 317 99 321
rect 0 316 99 317
rect 0 312 2 316
rect 96 312 99 316
rect 0 311 99 312
rect 0 307 2 311
rect 96 307 99 311
rect 0 306 99 307
rect 0 302 2 306
rect 96 302 99 306
rect 0 301 99 302
rect 0 297 2 301
rect 96 297 99 301
rect 0 296 99 297
rect 0 292 2 296
rect 96 292 99 296
rect 0 291 99 292
rect 0 287 2 291
rect 96 287 99 291
rect 0 286 99 287
rect 0 282 2 286
rect 96 282 99 286
rect 0 281 99 282
rect 0 277 2 281
rect 96 277 99 281
rect 0 276 99 277
rect 0 272 2 276
rect 96 272 99 276
rect 0 271 99 272
rect 0 267 2 271
rect 96 267 99 271
rect 0 266 99 267
rect 0 262 2 266
rect 96 262 99 266
rect 0 261 99 262
rect 0 257 7 261
rect 96 257 99 261
rect 0 256 99 257
rect 0 3 2 256
rect 6 252 8 256
rect 97 252 99 256
rect 6 251 99 252
rect 6 8 8 251
rect 102 248 140 329
rect 143 321 157 322
rect 143 316 157 317
rect 143 311 157 312
rect 143 306 157 307
rect 143 301 157 302
rect 143 296 157 297
rect 143 291 157 292
rect 143 286 157 287
rect 143 281 157 282
rect 143 276 157 277
rect 143 271 157 272
rect 143 266 157 267
rect 143 261 157 262
rect 143 256 157 257
rect 160 248 198 329
rect 201 322 204 326
rect 298 322 300 326
rect 201 321 300 322
rect 201 317 204 321
rect 298 317 300 321
rect 201 316 300 317
rect 201 312 204 316
rect 298 312 300 316
rect 201 311 300 312
rect 201 307 204 311
rect 298 307 300 311
rect 201 306 300 307
rect 201 302 204 306
rect 298 302 300 306
rect 201 301 300 302
rect 201 297 204 301
rect 298 297 300 301
rect 201 296 300 297
rect 201 292 204 296
rect 298 292 300 296
rect 201 291 300 292
rect 201 287 204 291
rect 298 287 300 291
rect 201 286 300 287
rect 201 282 204 286
rect 298 282 300 286
rect 201 281 300 282
rect 201 277 204 281
rect 298 277 300 281
rect 201 276 300 277
rect 201 272 204 276
rect 298 272 300 276
rect 201 271 300 272
rect 201 267 204 271
rect 298 267 300 271
rect 201 266 300 267
rect 201 262 204 266
rect 298 262 300 266
rect 201 261 300 262
rect 201 257 203 261
rect 292 257 300 261
rect 201 256 300 257
rect 201 252 203 256
rect 292 252 294 256
rect 201 251 294 252
rect 14 241 99 246
rect 14 237 19 241
rect 98 237 99 241
rect 14 233 99 237
rect 14 228 24 233
rect 14 29 19 228
rect 23 29 24 228
rect 28 229 39 233
rect 98 229 99 233
rect 28 227 99 229
rect 28 223 41 227
rect 95 223 99 227
rect 28 217 99 223
rect 28 43 32 217
rect 36 215 99 217
rect 36 196 39 215
rect 53 211 57 215
rect 96 211 99 215
rect 102 230 198 248
rect 102 208 142 230
rect 36 194 53 196
rect 36 175 39 194
rect 56 200 142 208
rect 157 208 198 230
rect 201 244 286 246
rect 201 235 202 244
rect 281 235 286 244
rect 201 233 286 235
rect 201 229 202 233
rect 261 229 277 233
rect 201 228 277 229
rect 201 227 272 228
rect 201 223 205 227
rect 259 223 272 227
rect 201 217 272 223
rect 201 215 264 217
rect 201 211 204 215
rect 243 211 247 215
rect 157 200 244 208
rect 120 196 180 200
rect 56 194 244 196
rect 120 190 180 194
rect 56 182 244 190
rect 261 196 264 215
rect 247 194 264 196
rect 53 175 57 179
rect 116 175 120 179
rect 36 167 120 175
rect 36 163 41 167
rect 36 161 120 163
rect 36 157 41 161
rect 36 149 120 157
rect 36 110 39 149
rect 53 145 57 149
rect 116 145 120 149
rect 123 142 177 182
rect 180 175 184 179
rect 243 175 247 179
rect 261 175 264 194
rect 180 167 264 175
rect 259 163 264 167
rect 180 161 264 163
rect 259 157 264 161
rect 180 149 264 157
rect 180 145 184 149
rect 243 145 247 149
rect 56 138 244 142
rect 56 134 142 138
rect 120 125 142 134
rect 56 120 142 125
rect 157 134 244 138
rect 157 125 180 134
rect 157 120 244 125
rect 56 117 244 120
rect 53 110 57 114
rect 116 110 120 114
rect 36 102 120 110
rect 36 98 41 102
rect 36 96 120 98
rect 36 92 41 96
rect 36 84 120 92
rect 36 45 39 84
rect 53 80 57 84
rect 116 80 120 84
rect 123 77 177 117
rect 180 110 184 114
rect 243 110 247 114
rect 261 110 264 149
rect 180 102 264 110
rect 259 98 264 102
rect 180 96 264 98
rect 259 92 264 96
rect 180 84 264 92
rect 180 80 184 84
rect 243 80 247 84
rect 56 70 244 77
rect 56 69 142 70
rect 120 60 142 69
rect 157 69 244 70
rect 56 52 142 60
rect 53 45 57 49
rect 96 45 99 49
rect 36 43 99 45
rect 28 37 99 43
rect 28 33 41 37
rect 95 33 99 37
rect 28 29 39 33
rect 98 29 99 33
rect 14 27 99 29
rect 14 23 19 27
rect 98 23 99 27
rect 14 22 99 23
rect 14 18 19 22
rect 98 18 99 22
rect 14 14 99 18
rect 102 28 142 52
rect 157 60 180 69
rect 157 52 244 60
rect 157 28 198 52
rect 6 7 99 8
rect 6 3 8 7
rect 92 3 99 7
rect 0 0 99 3
rect 102 0 198 28
rect 201 45 204 49
rect 243 45 247 49
rect 261 45 264 84
rect 201 43 264 45
rect 268 43 272 217
rect 201 37 272 43
rect 201 33 205 37
rect 259 33 272 37
rect 201 29 202 33
rect 261 29 272 33
rect 276 29 277 228
rect 281 29 286 233
rect 201 27 286 29
rect 201 23 202 27
rect 281 23 286 27
rect 201 22 286 23
rect 201 18 202 22
rect 281 18 286 22
rect 201 14 286 18
rect 292 8 294 251
rect 201 7 294 8
rect 201 3 203 7
rect 292 3 294 7
rect 298 3 300 256
rect 201 0 300 3
<< m2contact >>
rect 21 445 25 649
rect 36 638 120 642
rect 39 586 48 625
rect 52 621 116 625
rect 180 638 264 642
rect 184 621 248 625
rect 52 586 116 590
rect 39 522 48 561
rect 52 557 116 561
rect 143 606 157 610
rect 143 596 157 600
rect 184 586 248 590
rect 252 586 261 625
rect 184 557 248 561
rect 52 522 116 526
rect 39 457 48 496
rect 52 492 116 496
rect 143 542 157 546
rect 143 532 157 536
rect 184 522 248 526
rect 252 522 261 561
rect 184 492 248 496
rect 52 457 116 461
rect 143 477 157 481
rect 143 467 157 471
rect 184 457 248 461
rect 252 457 261 496
rect 275 445 279 649
rect 3 409 96 413
rect 3 399 96 403
rect 3 389 96 393
rect 3 379 96 383
rect 3 369 96 373
rect 3 359 96 363
rect 3 349 96 353
rect 143 409 157 413
rect 143 399 157 403
rect 143 389 157 393
rect 143 379 157 383
rect 143 369 157 373
rect 143 359 157 363
rect 143 349 157 353
rect 204 409 298 413
rect 204 399 298 403
rect 204 389 298 393
rect 204 379 298 383
rect 204 369 298 373
rect 204 359 298 363
rect 204 349 298 353
rect 2 317 96 321
rect 2 307 96 311
rect 2 297 96 301
rect 2 287 96 291
rect 2 277 96 281
rect 2 267 96 271
rect 7 257 96 261
rect 143 317 157 321
rect 143 307 157 311
rect 143 297 157 301
rect 143 287 157 291
rect 143 277 157 281
rect 143 267 157 271
rect 143 257 157 261
rect 204 317 298 321
rect 204 307 298 311
rect 204 297 298 301
rect 204 287 298 291
rect 204 277 298 281
rect 204 267 298 271
rect 203 257 292 261
rect 19 29 23 228
rect 39 196 53 215
rect 57 211 96 215
rect 39 175 53 194
rect 145 223 154 227
rect 145 215 154 219
rect 145 207 154 211
rect 204 211 243 215
rect 247 196 261 215
rect 57 175 116 179
rect 39 110 53 149
rect 57 145 116 149
rect 184 175 243 179
rect 247 175 261 194
rect 184 145 243 149
rect 145 127 154 131
rect 57 110 116 114
rect 39 45 53 84
rect 57 80 116 84
rect 184 110 243 114
rect 247 110 261 149
rect 184 80 243 84
rect 57 45 96 49
rect 39 29 98 33
rect 19 18 98 22
rect 145 63 154 67
rect 145 55 154 59
rect 145 47 154 51
rect 145 39 154 43
rect 145 31 154 35
rect 204 45 243 49
rect 247 45 261 84
rect 202 29 261 33
rect 272 29 276 228
rect 202 18 281 22
<< metal2 >>
rect 20 997 280 1000
rect 20 743 23 997
rect 277 743 280 997
rect 20 740 280 743
rect 0 649 300 670
rect 0 445 21 649
rect 25 642 275 649
rect 25 638 36 642
rect 120 638 180 642
rect 264 638 275 642
rect 25 625 275 638
rect 25 586 39 625
rect 48 621 52 625
rect 116 621 184 625
rect 248 621 252 625
rect 48 610 252 621
rect 48 606 143 610
rect 157 606 252 610
rect 48 600 252 606
rect 48 596 143 600
rect 157 596 252 600
rect 48 590 252 596
rect 48 586 52 590
rect 116 586 184 590
rect 248 586 252 590
rect 261 586 275 625
rect 25 561 275 586
rect 25 522 39 561
rect 48 557 52 561
rect 116 557 184 561
rect 248 557 252 561
rect 48 546 252 557
rect 48 542 143 546
rect 157 542 252 546
rect 48 536 252 542
rect 48 532 143 536
rect 157 532 252 536
rect 48 526 252 532
rect 48 522 52 526
rect 116 522 184 526
rect 248 522 252 526
rect 261 522 275 561
rect 25 496 275 522
rect 25 457 39 496
rect 48 492 52 496
rect 116 492 184 496
rect 248 492 252 496
rect 48 481 252 492
rect 48 477 143 481
rect 157 477 252 481
rect 48 471 252 477
rect 48 467 143 471
rect 157 467 252 471
rect 48 461 252 467
rect 48 457 52 461
rect 116 457 184 461
rect 248 457 252 461
rect 261 457 275 496
rect 25 445 275 457
rect 279 445 300 649
rect 0 440 300 445
rect 0 413 300 424
rect 0 409 3 413
rect 96 409 143 413
rect 157 409 204 413
rect 298 409 300 413
rect 0 403 300 409
rect 0 399 3 403
rect 96 399 143 403
rect 157 399 204 403
rect 298 399 300 403
rect 0 393 300 399
rect 0 389 3 393
rect 96 389 143 393
rect 157 389 204 393
rect 298 389 300 393
rect 0 383 300 389
rect 0 379 3 383
rect 96 379 143 383
rect 157 379 204 383
rect 298 379 300 383
rect 0 373 300 379
rect 0 369 3 373
rect 96 369 143 373
rect 157 369 204 373
rect 298 369 300 373
rect 0 363 300 369
rect 0 359 3 363
rect 96 359 143 363
rect 157 359 204 363
rect 298 359 300 363
rect 0 353 300 359
rect 0 349 3 353
rect 96 349 143 353
rect 157 349 204 353
rect 298 349 300 353
rect 0 344 300 349
rect 0 321 300 326
rect 0 317 2 321
rect 96 317 143 321
rect 157 317 204 321
rect 298 317 300 321
rect 0 311 300 317
rect 0 307 2 311
rect 96 307 143 311
rect 157 307 204 311
rect 298 307 300 311
rect 0 301 300 307
rect 0 297 2 301
rect 96 297 143 301
rect 157 297 204 301
rect 298 297 300 301
rect 0 291 300 297
rect 0 287 2 291
rect 96 287 143 291
rect 157 287 204 291
rect 298 287 300 291
rect 0 281 300 287
rect 0 277 2 281
rect 96 277 143 281
rect 157 277 204 281
rect 298 277 300 281
rect 0 271 300 277
rect 0 267 2 271
rect 96 267 143 271
rect 157 267 204 271
rect 298 267 300 271
rect 0 261 300 267
rect 0 257 7 261
rect 96 257 143 261
rect 157 257 203 261
rect 292 257 300 261
rect 0 246 300 257
rect 0 228 300 230
rect 0 29 19 228
rect 23 227 272 228
rect 23 223 145 227
rect 154 223 272 227
rect 23 219 272 223
rect 23 215 145 219
rect 154 215 272 219
rect 23 196 39 215
rect 53 211 57 215
rect 96 211 204 215
rect 243 211 247 215
rect 53 207 145 211
rect 154 207 247 211
rect 53 196 247 207
rect 261 196 272 215
rect 23 194 272 196
rect 23 175 39 194
rect 53 179 247 194
rect 53 175 57 179
rect 116 175 184 179
rect 243 175 247 179
rect 261 175 272 194
rect 23 149 272 175
rect 23 110 39 149
rect 53 145 57 149
rect 116 145 184 149
rect 243 145 247 149
rect 53 131 247 145
rect 53 127 145 131
rect 154 127 247 131
rect 53 114 247 127
rect 53 110 57 114
rect 116 110 184 114
rect 243 110 247 114
rect 261 110 272 149
rect 23 84 272 110
rect 23 45 39 84
rect 53 80 57 84
rect 116 80 184 84
rect 243 80 247 84
rect 53 67 247 80
rect 53 63 145 67
rect 154 63 247 67
rect 53 59 247 63
rect 53 55 145 59
rect 154 55 247 59
rect 53 51 247 55
rect 53 49 145 51
rect 53 45 57 49
rect 96 47 145 49
rect 154 49 247 51
rect 154 47 204 49
rect 96 45 204 47
rect 243 45 247 49
rect 261 45 272 84
rect 23 43 272 45
rect 23 39 145 43
rect 154 39 272 43
rect 23 35 272 39
rect 23 33 145 35
rect 23 29 39 33
rect 98 31 145 33
rect 154 33 272 35
rect 154 31 202 33
rect 98 29 202 31
rect 261 29 272 33
rect 276 29 300 228
rect 0 22 300 29
rect 0 18 19 22
rect 98 18 202 22
rect 281 18 300 22
rect 0 7 300 18
rect 0 0 98 7
rect 202 0 300 7
<< pad >>
rect 23 743 277 997
<< m1p >>
rect 102 0 198 4
<< m3p >>
rect 144 868 167 891
<< labels >>
rlabel m3p 155 879 155 879 1 YPAD
rlabel m1p 150 0 150 0 1 POWER
<< end >>
