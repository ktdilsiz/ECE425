magic
tech scmos
timestamp 1485568973
<< nwell >>
rect -6 40 26 96
<< ntransistor >>
rect 5 7 7 23
rect 13 7 15 23
<< ptransistor >>
rect 5 51 7 83
rect 10 51 12 83
<< ndiffusion >>
rect 0 22 5 23
rect 4 8 5 22
rect 0 7 5 8
rect 7 22 13 23
rect 7 8 8 22
rect 12 8 13 22
rect 7 7 13 8
rect 15 22 20 23
rect 15 8 16 22
rect 15 7 20 8
<< pdiffusion >>
rect 0 81 5 83
rect 4 52 5 81
rect 0 51 5 52
rect 7 51 10 83
rect 12 81 17 83
rect 12 52 13 81
rect 12 51 17 52
<< ndcontact >>
rect 0 8 4 22
rect 8 8 12 22
rect 16 8 20 22
<< pdcontact >>
rect 0 52 4 81
rect 13 52 17 81
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
<< polysilicon >>
rect 5 83 7 85
rect 10 83 12 85
rect 5 23 7 51
rect 10 44 12 51
rect 10 42 15 44
rect 13 23 15 42
rect 5 5 7 7
rect 13 5 15 7
<< polycontact >>
rect 1 43 5 47
rect 15 26 19 30
<< metal1 >>
rect -2 92 22 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 22 92
rect -2 86 22 88
rect 0 81 4 86
rect 0 51 4 52
rect 13 81 17 83
rect 13 37 17 52
rect 12 33 17 37
rect 0 22 4 23
rect 0 4 4 8
rect 8 22 12 33
rect 8 7 12 8
rect 16 22 20 23
rect 16 4 20 8
rect -2 2 22 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 22 2
rect -2 -4 22 -2
<< m2contact >>
rect 0 43 1 47
rect 1 43 4 47
rect 8 33 12 37
rect 16 26 19 30
rect 19 26 20 30
<< labels >>
rlabel metal1 -1 0 -1 0 2 Gnd!
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel m2contact 1 45 1 45 1 a
rlabel m2contact 10 35 10 35 1 y
rlabel m2contact 18 28 18 28 1 b
<< end >>
