magic
tech scmos
timestamp 1484532969
<< nwell >>
rect -6 40 34 96
<< ntransistor >>
rect 5 7 7 34
rect 21 7 23 34
<< ptransistor >>
rect 5 46 7 83
rect 21 46 23 83
<< ndiffusion >>
rect 0 32 5 34
rect 4 8 5 32
rect 0 7 5 8
rect 7 32 12 34
rect 7 8 8 32
rect 7 7 12 8
rect 16 32 21 34
rect 20 8 21 32
rect 16 7 21 8
rect 23 32 28 34
rect 23 8 24 32
rect 23 7 28 8
<< pdiffusion >>
rect 0 81 5 83
rect 4 47 5 81
rect 0 46 5 47
rect 7 81 12 83
rect 7 47 8 81
rect 7 46 12 47
rect 16 81 21 83
rect 20 47 21 81
rect 16 46 21 47
rect 23 81 28 83
rect 23 47 24 81
rect 23 46 28 47
<< ndcontact >>
rect 0 8 4 32
rect 8 8 12 32
rect 16 8 20 32
rect 24 8 28 32
<< pdcontact >>
rect 0 47 4 81
rect 8 47 12 81
rect 16 47 20 81
rect 24 47 28 81
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
<< polysilicon >>
rect 5 83 7 85
rect 21 83 23 85
rect 5 34 7 46
rect 21 41 23 46
rect 17 39 23 41
rect 21 34 23 39
rect 5 5 7 7
rect 21 5 23 7
<< polycontact >>
rect 1 38 5 42
rect 13 38 17 42
<< metal1 >>
rect -2 92 30 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 30 92
rect -2 86 30 88
rect 0 81 4 86
rect 0 46 4 47
rect 8 81 12 83
rect 8 42 12 47
rect 16 81 20 86
rect 16 46 20 47
rect 24 81 28 83
rect 24 42 28 47
rect 12 38 13 42
rect 0 32 4 34
rect 0 4 4 8
rect 8 32 12 38
rect 8 7 12 8
rect 16 32 20 34
rect 16 4 20 8
rect 24 32 28 38
rect 24 7 28 8
rect -2 2 30 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 30 2
rect -2 -4 30 -2
<< m2contact >>
rect 0 38 1 42
rect 1 38 4 42
rect 8 38 12 42
rect 24 38 28 42
<< labels >>
rlabel m2contact 1 40 1 40 1 s
rlabel m2contact 10 40 10 40 1 sb_out
rlabel m2contact 26 40 26 40 1 s_out
rlabel metal1 -1 0 -1 0 3 Gnd!
rlabel metal1 -1 90 -1 90 3 Vdd!
<< end >>
