magic
tech scmos
timestamp 1487715524
<< nwell >>
rect -4 40 36 96
<< ntransistor >>
rect 7 7 9 11
rect 12 7 14 11
rect 20 7 22 11
<< ptransistor >>
rect 7 79 9 83
rect 15 79 17 83
rect 23 79 25 83
<< ndiffusion >>
rect 6 7 7 11
rect 9 7 12 11
rect 14 7 15 11
rect 19 7 20 11
rect 22 7 23 11
<< pdiffusion >>
rect 6 79 7 83
rect 9 79 10 83
rect 14 79 15 83
rect 17 79 18 83
rect 22 79 23 83
rect 25 79 26 83
<< ndcontact >>
rect 2 7 6 11
rect 15 7 19 11
rect 23 7 27 11
<< pdcontact >>
rect 2 79 6 83
rect 10 79 14 83
rect 18 79 22 83
rect 26 79 30 83
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 88 6 92
rect 10 88 14 92
rect 18 88 22 92
rect 26 88 30 92
<< polysilicon >>
rect 7 83 9 85
rect 15 83 17 85
rect 23 83 25 85
rect 7 62 9 79
rect 15 62 17 79
rect 23 78 25 79
rect 2 60 9 62
rect 12 60 17 62
rect 20 76 25 78
rect 2 37 4 60
rect 12 37 14 60
rect 20 37 22 76
rect 26 33 30 37
rect 2 24 4 33
rect 2 22 9 24
rect 7 11 9 22
rect 12 11 14 33
rect 20 11 22 33
rect 7 5 9 7
rect 12 5 14 7
rect 20 5 22 7
<< polycontact >>
rect 2 33 6 37
rect 10 33 14 37
rect 18 33 22 37
<< metal1 >>
rect 0 92 32 94
rect 0 88 2 92
rect 6 88 10 92
rect 14 88 18 92
rect 22 88 26 92
rect 30 88 32 92
rect 0 86 32 88
rect 10 83 14 86
rect 2 75 6 79
rect 18 75 22 79
rect 2 71 22 75
rect 26 37 30 79
rect 26 21 30 33
rect 15 17 30 21
rect 15 11 19 17
rect 2 4 6 7
rect 23 4 27 7
rect 0 2 32 4
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 32 2
rect 0 -4 32 -2
<< m2contact >>
rect 2 33 6 37
rect 10 33 14 37
rect 18 33 22 37
rect 26 33 30 37
<< labels >>
rlabel m2contact 4 35 4 35 1 a
rlabel m2contact 12 35 12 35 1 b
rlabel m2contact 20 35 20 35 1 c
rlabel metal1 1 0 1 0 2 Gnd!
rlabel metal1 1 90 1 90 3 Vdd!
rlabel m2contact 28 35 28 35 1 y
<< end >>
