magic
tech scmos
timestamp 1484435125
<< nwell >>
rect -6 40 50 96
<< ntransistor >>
rect 10 7 12 13
rect 15 7 17 13
rect 23 7 25 13
rect 28 7 30 13
rect 36 7 38 14
<< ptransistor >>
rect 10 74 12 83
rect 15 74 17 83
rect 23 74 25 83
rect 28 74 30 83
rect 36 73 38 83
<< ndiffusion >>
rect 31 13 36 14
rect 5 12 10 13
rect 9 8 10 12
rect 5 7 10 8
rect 12 7 15 13
rect 17 12 23 13
rect 17 8 18 12
rect 22 8 23 12
rect 17 7 23 8
rect 25 7 28 13
rect 30 12 36 13
rect 30 8 31 12
rect 35 8 36 12
rect 30 7 36 8
rect 38 12 43 14
rect 38 8 39 12
rect 38 7 43 8
<< pdiffusion >>
rect 9 74 10 83
rect 12 74 15 83
rect 17 74 18 83
rect 22 74 23 83
rect 25 74 28 83
rect 30 82 36 83
rect 30 74 31 82
rect 35 73 36 82
rect 38 82 43 83
rect 38 73 39 82
<< ndcontact >>
rect 5 8 9 12
rect 18 8 22 12
rect 31 8 35 12
rect 39 8 43 12
<< pdcontact >>
rect 5 74 9 83
rect 18 74 22 83
rect 31 73 35 82
rect 39 73 43 82
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
rect 40 -2 44 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
rect 32 88 36 92
rect 40 88 44 92
<< polysilicon >>
rect 10 83 12 85
rect 15 83 17 85
rect 23 83 25 85
rect 28 83 30 85
rect 36 83 38 85
rect 10 65 12 74
rect 2 63 12 65
rect 2 50 4 63
rect 15 60 17 74
rect 9 58 17 60
rect 9 50 11 58
rect 23 55 25 74
rect 18 53 25 55
rect 28 49 30 74
rect 2 16 4 46
rect 18 42 20 49
rect 15 40 20 42
rect 2 14 12 16
rect 10 13 12 14
rect 15 13 17 40
rect 27 33 29 45
rect 36 41 38 73
rect 37 37 38 41
rect 27 31 31 33
rect 23 13 25 23
rect 29 17 31 31
rect 28 15 31 17
rect 28 13 30 15
rect 36 14 38 37
rect 10 5 12 7
rect 15 5 17 7
rect 23 5 25 7
rect 28 5 30 7
rect 36 5 38 7
<< polycontact >>
rect 0 46 4 50
rect 8 46 12 50
rect 18 49 22 53
rect 26 45 30 49
rect 33 37 37 41
rect 21 23 25 27
<< metal1 >>
rect -2 92 46 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 32 92
rect 36 88 40 92
rect 44 88 46 92
rect -2 86 46 88
rect 5 83 9 86
rect 18 69 22 74
rect 31 82 35 86
rect 39 82 43 83
rect 20 65 22 69
rect 18 55 24 59
rect 18 53 22 55
rect 39 50 43 73
rect 8 27 12 46
rect 30 45 32 48
rect 26 44 32 45
rect 39 46 44 50
rect 40 42 44 46
rect 31 37 33 41
rect 31 35 35 37
rect 20 32 35 35
rect 20 31 27 32
rect 31 31 35 32
rect 40 31 44 38
rect 39 27 44 31
rect 8 23 21 27
rect 20 15 22 19
rect 5 12 9 13
rect 5 4 9 8
rect 18 12 22 15
rect 18 7 22 8
rect 31 12 35 14
rect 31 4 35 8
rect 39 12 43 27
rect 39 7 43 8
rect -2 2 46 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 40 2
rect 44 -2 46 2
rect -2 -4 46 -2
<< m2contact >>
rect 16 65 20 69
rect 24 55 28 59
rect 0 46 4 50
rect 8 46 12 50
rect 32 44 36 48
rect 40 38 44 42
rect 16 31 20 35
rect 16 15 20 19
<< metal2 >>
rect 16 35 20 65
rect 16 19 20 31
<< labels >>
rlabel metal1 -1 0 -1 0 2 Gnd!
rlabel m2contact 42 40 42 40 1 y
rlabel m2contact 34 46 34 46 1 d0
rlabel m2contact 26 57 26 57 1 s
rlabel m2contact 10 48 10 48 1 sb
rlabel m2contact 2 48 2 48 1 d1
rlabel metal1 -1 90 -1 90 3 Vdd!
<< end >>
