magic
tech scmos
timestamp 1484455428
<< nwell >>
rect -6 40 42 96
<< ntransistor >>
rect 5 7 7 16
rect 21 7 23 25
rect 29 7 31 25
<< ptransistor >>
rect 5 65 7 83
rect 21 47 23 83
rect 29 47 31 83
<< ndiffusion >>
rect 16 23 21 25
rect 4 7 5 16
rect 7 7 8 16
rect 20 9 21 23
rect 16 7 21 9
rect 23 23 29 25
rect 23 9 24 23
rect 28 9 29 23
rect 23 7 29 9
rect 31 23 36 25
rect 31 9 32 23
rect 31 7 36 9
<< pdiffusion >>
rect 0 81 5 83
rect 4 67 5 81
rect 0 65 5 67
rect 7 81 12 83
rect 7 67 8 81
rect 7 65 12 67
rect 16 82 21 83
rect 20 49 21 82
rect 16 47 21 49
rect 23 82 29 83
rect 23 48 24 82
rect 28 48 29 82
rect 23 47 29 48
rect 31 82 36 83
rect 31 49 32 82
rect 31 47 36 49
<< ndcontact >>
rect 0 7 4 16
rect 8 7 12 16
rect 16 9 20 23
rect 24 9 28 23
rect 32 9 36 23
<< pdcontact >>
rect 0 67 4 81
rect 8 67 12 81
rect 16 49 20 82
rect 24 48 28 82
rect 32 49 36 82
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
rect 32 88 36 92
<< polysilicon >>
rect 5 83 7 85
rect 21 83 23 85
rect 29 83 31 85
rect 5 59 7 65
rect 1 30 3 58
rect 21 30 23 47
rect 29 42 31 47
rect 1 28 23 30
rect 5 16 7 28
rect 21 25 23 28
rect 29 25 31 38
rect 5 5 7 7
rect 21 5 23 7
rect 29 5 31 7
<< polycontact >>
rect 1 58 5 62
rect 28 38 32 42
<< metal1 >>
rect -2 92 38 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 32 92
rect 36 88 38 92
rect -2 86 38 88
rect 0 81 4 86
rect 0 65 4 67
rect 8 81 12 83
rect 8 42 12 67
rect 16 82 20 83
rect 24 82 28 86
rect 24 47 28 48
rect 32 82 36 83
rect 8 38 28 42
rect 8 16 12 38
rect 16 7 20 9
rect 24 23 28 25
rect 0 4 4 7
rect 24 4 28 9
rect 32 7 36 9
rect -2 2 38 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 38 2
rect -2 -4 38 -2
<< m2contact >>
rect 0 58 1 62
rect 1 58 4 62
rect 16 49 20 51
rect 16 47 20 49
rect 32 49 36 51
rect 32 47 36 49
rect 16 23 20 25
rect 16 21 20 23
rect 32 23 36 25
rect 32 21 36 23
<< metal2 >>
rect 16 25 20 47
rect 32 25 36 47
<< labels >>
rlabel m2contact 2 60 2 60 1 ph
rlabel m2contact 18 23 18 23 1 phb
rlabel m2contact 34 23 34 23 1 phbuf
rlabel metal1 -1 -1 -1 0 2 Gnd!
rlabel metal1 -1 90 -1 90 3 Vdd!
<< end >>
