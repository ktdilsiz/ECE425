magic
tech scmos
timestamp 1488311641
<< nwell >>
rect -8 48 16 105
<< psubstratepcontact >>
rect -2 -2 2 2
rect 6 -2 10 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 6 98 10 102
<< metal1 >>
rect -2 102 10 103
rect 2 98 6 102
rect -2 97 10 98
rect -2 2 10 3
rect 2 -2 6 2
rect -2 -3 10 -2
<< labels >>
flabel metal1 4 100 4 100 4 FreeSans 26 0 0 0 vdd
flabel metal1 4 0 4 0 4 FreeSans 26 0 0 0 gnd
<< end >>
