magic
tech scmos
timestamp 1484539914
<< metal1 >>
rect -153 338 1131 340
rect -89 334 1111 338
rect 1130 334 1131 338
rect -153 332 1131 334
rect 2724 338 2788 340
rect 2724 332 2788 334
rect -243 326 367 328
rect -179 322 367 326
rect -243 320 367 322
rect 2634 326 2698 328
rect 2634 320 2698 322
rect -243 203 6 205
rect -179 199 172 203
rect -243 197 6 199
rect -153 113 6 115
rect -89 109 172 113
rect -153 107 6 109
rect -243 92 6 94
rect -179 88 172 92
rect -243 86 6 88
rect 359 4 367 320
rect 2634 203 2698 205
rect 2634 197 2698 199
rect 2724 113 2788 115
rect 2724 107 2788 109
rect 1047 92 2698 94
rect 1066 88 2634 92
rect 1047 86 2698 88
rect -153 2 6 4
rect 359 2 1067 4
rect -89 -2 172 2
rect 359 -2 1047 2
rect 1066 -2 1067 2
rect -153 -4 6 -2
rect 359 -4 1067 -2
rect 1111 2 2788 4
rect 1130 -2 2724 2
rect 1111 -4 2788 -2
rect 4 -30 744 -26
rect 772 -30 1808 -26
rect 740 -38 960 -34
rect 1534 -38 2048 -34
rect 588 -46 664 -42
rect 716 -46 1960 -42
rect 700 -54 1992 -50
rect 228 -62 476 -58
rect 700 -62 760 -58
rect 1502 -62 2216 -58
rect 220 -70 460 -66
rect 724 -70 792 -66
rect 1574 -70 2240 -66
rect 212 -78 444 -74
rect 732 -78 1602 -74
rect 204 -86 428 -82
rect 740 -86 1594 -82
rect 1654 -86 2480 -82
rect 196 -94 412 -90
rect 748 -94 1538 -90
rect 1590 -94 2512 -90
rect 188 -102 396 -98
rect 428 -102 648 -98
rect 756 -102 1618 -98
rect 244 -110 640 -106
rect 676 -110 1632 -106
rect 60 -118 624 -114
rect 692 -118 1600 -114
<< m2contact >>
rect -153 334 -89 338
rect 1111 334 1130 338
rect 2724 334 2788 338
rect -243 322 -179 326
rect 2634 322 2698 326
rect -243 199 -179 203
rect -153 109 -89 113
rect -243 88 -179 92
rect 2634 199 2698 203
rect 2724 109 2788 113
rect 1047 88 1066 92
rect 2634 88 2698 92
rect -153 -2 -89 2
rect 1047 -2 1066 2
rect 1111 -2 1130 2
rect 2724 -2 2788 2
rect 0 -30 4 -26
rect 744 -30 748 -26
rect 768 -30 772 -26
rect 1808 -30 1812 -26
rect 736 -38 740 -34
rect 960 -38 964 -34
rect 1530 -38 1534 -34
rect 2048 -38 2052 -34
rect 584 -46 588 -42
rect 664 -46 668 -42
rect 712 -46 716 -42
rect 1960 -46 1964 -42
rect 696 -54 700 -50
rect 1992 -54 1996 -50
rect 224 -62 228 -58
rect 476 -62 480 -58
rect 696 -62 700 -58
rect 760 -62 764 -58
rect 1498 -62 1502 -58
rect 2216 -62 2220 -58
rect 216 -70 220 -66
rect 460 -70 464 -66
rect 720 -70 724 -66
rect 792 -70 796 -66
rect 1570 -70 1574 -66
rect 2240 -70 2244 -66
rect 208 -78 212 -74
rect 444 -78 448 -74
rect 728 -78 732 -74
rect 1602 -78 1606 -74
rect 200 -86 204 -82
rect 428 -86 432 -82
rect 736 -86 740 -82
rect 1594 -86 1598 -82
rect 1650 -86 1654 -82
rect 2480 -86 2484 -82
rect 192 -94 196 -90
rect 412 -94 416 -90
rect 744 -94 748 -90
rect 1538 -94 1542 -90
rect 1586 -94 1590 -90
rect 2512 -94 2516 -90
rect 184 -102 188 -98
rect 396 -102 400 -98
rect 424 -102 428 -98
rect 648 -102 652 -98
rect 752 -102 756 -98
rect 1618 -102 1622 -98
rect 240 -110 244 -106
rect 640 -110 644 -106
rect 672 -110 676 -106
rect 1632 -110 1636 -106
rect 56 -118 60 -114
rect 624 -118 628 -114
rect 688 -118 692 -114
rect 1600 -118 1604 -114
<< metal2 >>
rect -243 326 -179 355
rect -243 203 -179 322
rect -243 92 -179 199
rect -243 -172 -179 88
rect -153 338 -89 368
rect -153 113 -89 334
rect 1111 338 1131 346
rect 1130 334 1131 338
rect -33 171 -27 172
rect -33 167 -32 171
rect -28 167 -27 171
rect 135 171 141 172
rect 135 167 136 171
rect 140 167 141 171
rect 303 171 309 172
rect 303 167 304 171
rect 308 167 309 171
rect -33 166 -27 167
rect 0 153 4 167
rect 135 166 141 167
rect -41 152 -35 153
rect -41 148 -40 152
rect -36 148 -35 152
rect -41 147 -35 148
rect -17 152 -11 153
rect -1 152 5 153
rect -17 148 -16 152
rect -12 148 -11 152
rect -8 148 0 152
rect 4 148 5 152
rect -17 147 -11 148
rect -1 147 5 148
rect -25 122 -19 123
rect -25 118 -24 122
rect -20 118 -19 122
rect -25 117 -19 118
rect -153 2 -89 109
rect 0 54 4 147
rect 8 132 12 157
rect 7 131 13 132
rect 7 127 8 131
rect 12 127 13 131
rect 7 126 13 127
rect 24 123 28 157
rect 23 122 29 123
rect 23 118 24 122
rect 28 118 29 122
rect 23 117 29 118
rect 8 23 12 47
rect 24 44 28 117
rect 136 30 140 166
rect 159 162 165 163
rect 159 158 160 162
rect 164 158 165 162
rect 159 157 165 158
rect 160 150 164 157
rect 168 153 172 167
rect 303 166 309 167
rect 167 152 173 153
rect 167 148 168 152
rect 172 148 173 152
rect 167 147 173 148
rect 168 54 172 147
rect 176 143 180 157
rect 175 142 181 143
rect 175 138 176 142
rect 180 138 181 142
rect 175 137 181 138
rect 192 123 196 157
rect 191 122 197 123
rect 191 118 192 122
rect 196 118 197 122
rect 191 117 197 118
rect 159 52 165 53
rect 159 48 160 52
rect 164 48 165 52
rect 159 47 165 48
rect 160 39 164 47
rect 176 43 180 47
rect 192 44 196 117
rect 175 42 181 43
rect 175 38 176 42
rect 180 38 181 42
rect 175 37 181 38
rect 304 30 308 166
rect 491 162 497 163
rect 491 158 492 162
rect 496 158 497 162
rect 491 157 497 158
rect 328 152 334 153
rect 328 148 329 152
rect 333 148 334 152
rect 328 147 334 148
rect 328 42 334 43
rect 328 38 329 42
rect 333 38 334 42
rect 328 37 334 38
rect 7 22 13 23
rect 7 18 8 22
rect 12 18 13 22
rect 7 17 13 18
rect -153 -172 -89 -2
rect 0 -142 4 -30
rect 56 -142 60 -118
rect 184 -142 188 -102
rect 192 -142 196 -94
rect 200 -142 204 -86
rect 208 -142 212 -78
rect 216 -142 220 -70
rect 224 -142 228 -62
rect 396 -98 400 25
rect 412 -90 416 25
rect 428 -82 432 25
rect 444 -74 448 25
rect 460 -66 464 25
rect 476 -58 480 25
rect 492 23 496 157
rect 523 152 529 153
rect 523 148 524 152
rect 528 148 529 152
rect 523 147 529 148
rect 507 52 513 53
rect 507 48 508 52
rect 512 48 513 52
rect 507 47 513 48
rect 508 23 512 47
rect 524 23 528 147
rect 831 142 837 143
rect 831 138 832 142
rect 836 138 837 142
rect 831 137 837 138
rect 807 132 813 133
rect 807 128 808 132
rect 812 128 813 132
rect 807 127 813 128
rect 575 72 581 73
rect 575 68 576 72
rect 580 68 581 72
rect 575 67 581 68
rect 539 42 545 43
rect 539 38 540 42
rect 544 38 545 42
rect 539 37 545 38
rect 540 23 544 37
rect 576 23 580 67
rect 591 62 597 63
rect 591 58 592 62
rect 596 58 597 62
rect 591 57 597 58
rect 592 23 596 57
rect 615 52 621 53
rect 615 48 616 52
rect 620 48 621 52
rect 615 47 621 48
rect 599 42 605 43
rect 599 38 600 42
rect 604 38 605 42
rect 599 37 605 38
rect 600 23 604 37
rect 616 23 620 47
rect 240 -142 244 -110
rect 424 -142 428 -102
rect 584 -142 588 -46
rect 624 -114 628 25
rect 640 -106 644 25
rect 648 -98 652 25
rect 664 -42 668 25
rect 672 -106 676 25
rect 688 -114 692 25
rect 696 -50 700 25
rect 712 -42 716 25
rect 696 -142 700 -62
rect 720 -66 724 25
rect 736 -34 740 25
rect 744 -26 748 25
rect 760 -58 764 25
rect 768 -26 772 25
rect 784 -57 788 25
rect 792 -17 796 25
rect 808 23 812 127
rect 816 23 820 25
rect 832 23 836 137
rect 1047 92 1067 100
rect 1066 88 1067 92
rect 839 32 845 33
rect 839 28 840 32
rect 844 28 845 32
rect 839 27 845 28
rect 840 23 844 27
rect 815 22 821 23
rect 815 18 816 22
rect 820 18 821 22
rect 815 17 821 18
rect 1047 2 1067 88
rect 1066 -2 1067 2
rect 1047 -10 1067 -2
rect 1111 2 1131 334
rect 2634 326 2698 355
rect 2634 203 2698 322
rect 2634 92 2698 199
rect 1545 72 1551 73
rect 1545 68 1546 72
rect 1550 68 1551 72
rect 1545 67 1551 68
rect 1513 52 1519 53
rect 1513 48 1514 52
rect 1518 48 1519 52
rect 1513 47 1519 48
rect 1130 -2 1131 2
rect 1111 -11 1131 -2
rect 791 -18 797 -17
rect 791 -22 792 -18
rect 796 -22 797 -18
rect 791 -23 797 -22
rect 783 -58 789 -57
rect 783 -62 784 -58
rect 788 -62 789 -58
rect 783 -63 789 -62
rect 728 -142 732 -78
rect 736 -142 740 -86
rect 744 -142 748 -94
rect 752 -142 756 -102
rect 792 -142 796 -70
rect 960 -142 964 -38
rect 1498 -58 1502 47
rect 1506 43 1510 46
rect 1514 44 1518 47
rect 1505 42 1511 43
rect 1505 38 1506 42
rect 1510 38 1511 42
rect 1505 37 1511 38
rect 1530 -34 1534 50
rect 1546 43 1550 67
rect 1553 62 1559 63
rect 1553 58 1554 62
rect 1558 58 1559 62
rect 1553 57 1559 58
rect 1554 43 1558 57
rect 1538 -90 1542 -8
rect 1570 -66 1574 -8
rect 1586 -90 1590 -8
rect 1594 -82 1598 -8
rect 1602 -74 1606 -8
rect 1618 -98 1622 -8
rect 1650 -82 1654 -8
rect 1600 -142 1604 -118
rect 1632 -142 1636 -110
rect 1808 -142 1812 -30
rect 1960 -142 1964 -46
rect 1992 -142 1996 -54
rect 2048 -142 2052 -38
rect 2216 -142 2220 -62
rect 2240 -142 2244 -70
rect 2480 -142 2484 -86
rect 2512 -142 2516 -94
rect 2634 -172 2698 88
rect 2724 338 2788 368
rect 2724 113 2788 334
rect 2724 2 2788 109
rect 2724 -172 2788 -2
<< m3contact >>
rect -32 167 -28 171
rect 136 167 140 171
rect 304 167 308 171
rect -40 148 -36 152
rect -16 148 -12 152
rect 0 148 4 152
rect -24 118 -20 122
rect 8 127 12 131
rect 24 118 28 122
rect 160 158 164 162
rect 168 148 172 152
rect 176 138 180 142
rect 192 118 196 122
rect 160 48 164 52
rect 176 38 180 42
rect 492 158 496 162
rect 329 148 333 152
rect 329 38 333 42
rect 8 18 12 22
rect 524 148 528 152
rect 508 48 512 52
rect 832 138 836 142
rect 808 128 812 132
rect 576 68 580 72
rect 540 38 544 42
rect 592 58 596 62
rect 616 48 620 52
rect 600 38 604 42
rect 840 28 844 32
rect 816 18 820 22
rect 1546 68 1550 72
rect 1514 48 1518 52
rect 792 -22 796 -18
rect 784 -62 788 -58
rect 1506 38 1510 42
rect 1554 58 1558 62
<< metal3 >>
rect -33 171 309 172
rect -33 167 -32 171
rect -28 167 136 171
rect 140 167 304 171
rect 308 167 309 171
rect -33 166 309 167
rect 159 162 497 163
rect 159 158 160 162
rect 164 158 492 162
rect 496 158 497 162
rect 159 157 497 158
rect -41 152 -11 153
rect -41 148 -40 152
rect -36 148 -16 152
rect -12 148 -11 152
rect -41 147 -11 148
rect -1 152 173 153
rect -1 148 0 152
rect 4 148 168 152
rect 172 148 173 152
rect -1 147 173 148
rect 328 152 529 153
rect 328 148 329 152
rect 333 148 524 152
rect 528 148 529 152
rect 328 147 529 148
rect 175 142 837 143
rect 175 138 176 142
rect 180 138 832 142
rect 836 138 837 142
rect 175 137 837 138
rect 7 132 813 133
rect 7 131 808 132
rect 7 127 8 131
rect 12 128 808 131
rect 812 128 813 132
rect 12 127 813 128
rect 7 126 13 127
rect -25 122 197 123
rect -25 118 -24 122
rect -20 118 24 122
rect 28 118 192 122
rect 196 118 197 122
rect -25 117 197 118
rect 575 72 1551 73
rect 575 68 576 72
rect 580 68 1546 72
rect 1550 68 1551 72
rect 575 67 1551 68
rect 591 62 1559 63
rect 591 58 592 62
rect 596 58 1554 62
rect 1558 58 1559 62
rect 591 57 1559 58
rect 159 52 513 53
rect 159 48 160 52
rect 164 48 508 52
rect 512 48 513 52
rect 159 47 513 48
rect 615 52 1519 53
rect 615 48 616 52
rect 620 48 1514 52
rect 1518 48 1519 52
rect 615 47 1519 48
rect 175 42 181 43
rect 175 38 176 42
rect 180 38 181 42
rect 175 33 181 38
rect 328 42 545 43
rect 328 38 329 42
rect 333 38 540 42
rect 544 38 545 42
rect 328 37 545 38
rect 599 42 1511 43
rect 599 38 600 42
rect 604 38 1506 42
rect 1510 38 1511 42
rect 599 37 1511 38
rect 175 32 845 33
rect 175 28 840 32
rect 844 28 845 32
rect 175 27 845 28
rect 7 22 821 23
rect 7 18 8 22
rect 12 18 816 22
rect 820 18 821 22
rect 7 17 821 18
rect -13 -18 797 -17
rect -13 -22 792 -18
rect 796 -22 797 -18
rect -13 -23 797 -22
rect -13 -58 789 -57
rect -13 -62 784 -58
rect 788 -62 789 -58
rect -13 -63 789 -62
use inv_1x  inv_1x_0
timestamp 1484418501
transform 1 0 -16 0 1 111
box -6 -4 18 96
use flopr_c_1x  flopr_c_1x_0
timestamp 1484536911
transform 1 0 -24 0 1 111
box 18 -4 194 96
use flopr_c_1x  flopr_c_1x_1
timestamp 1484536911
transform 1 0 144 0 1 111
box 18 -4 194 96
use flopr_c_1x  flopr_c_1x_2
timestamp 1484536911
transform 1 0 -24 0 1 0
box 18 -4 194 96
use flopr_c_1x  flopr_c_1x_3
timestamp 1484536911
transform 1 0 144 0 1 0
box 18 -4 194 96
use controller_pla  controller_pla_0
timestamp 1484539528
transform 1 0 361 0 1 0
box -6 -8 497 340
use a2o1_1x  a2o1_1x_0
timestamp 1484539914
transform 1 0 1498 0 1 0
box -6 -4 42 96
use aludec  aludec_0
timestamp 1484539914
transform 1 0 1538 0 1 0
box -6 -12 130 112
<< end >>
