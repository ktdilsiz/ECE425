alu_decoder_testbench.sv                                                                            0000644 �    Asz0000145 00000002617 13055345410 013661  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   `timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/28/2017 01:59:08 PM
// Design Name: 
// Module Name: alu_decoder_testbench
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module alu_decoder_testbench();

logic [1:0] alu_op;
logic [5:0] funct;
logic [6:0] op;
logic clk;
    alu_ctl DUV_aluctl(.alu_op(alu_op), .funct(funct), .op(op));
    
  always
     begin
	clk = 0;
	#10 clk = 1;
	#10 ;
end

    initial begin
    
        alu_op=00;
        @(posedge clk);
        alu_op=00;
        @(posedge clk);
        alu_op=01;
        @(posedge clk);
        alu_op=10;
        funct = 6'h20;
        @(posedge clk);
        alu_op=10;
        funct = 6'h20;
        @(posedge clk);
        alu_op=10;
        funct = 6'h22;
        @(posedge clk);
        alu_op=10;
        funct = 6'h24;
        @(posedge clk);
        alu_op=10;
        funct = 6'h25;
        @(posedge clk);
        alu_op=10;
        funct = 6'h26;
        @(posedge clk);
        alu_op=10;
        funct = 6'h27;
        @(posedge clk);
        alu_op=10;
        funct = 6'h2b;  
        end                              

endmodule
                                                                                                                 alu_ctl.nofill.v                                                                                    0000644 �    Asz0000145 00000004451 13055352430 012074  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   //
// Milkyway Hierarchical Verilog Dump:
// Generated on 02/28/2017 at 14:52:56
// Design Generated by Consolidated Verilog Reader
// File produced by Consolidated Verilog Writer
// Library Name :alu_ctl_LIB
// Cell Name    :alu_ctl
// Hierarchy delimiter:'/'
// Write Command : write_verilog alu_ctl.pnr.v
//


module alu_ctl (funct , alu_op , op );
input  [5:0] funct ;
input  [1:0] alu_op ;
output [6:0] op ;



INVX2 U10 (.A ( funct[1] ) , .Y ( n7 ) ) ;
INVX2 U9 (.A ( funct[2] ) , .Y ( n6 ) ) ;
INVX2 U8 (.A ( n17 ) , .Y ( n5 ) ) ;
INVX2 U7 (.A ( n15 ) , .Y ( n4 ) ) ;
INVX2 U6 (.A ( n22 ) , .Y ( op[1] ) ) ;
INVX2 U5 (.A ( alu_op[1] ) , .Y ( n2 ) ) ;
INVX2 U4 (.A ( op[2] ) , .Y ( n1 ) ) ;
AND2X2 U3 (.A ( funct[1] ) , .B ( funct[3] ) , .Y ( n24 ) ) ;
OAI21X1 U18 (.A ( n5 ) , .B ( n15 ) , .C ( n16 ) , .Y ( op[4] ) ) ;
XOR2X1 U17 (.A ( funct[2] ) , .B ( funct[1] ) , .Y ( n13 ) ) ;
OAI21X1 U16 (.A ( funct[0] ) , .B ( n13 ) , .C ( n14 ) , .Y ( n12 ) ) ;
NAND2X1 U15 (.A ( n11 ) , .B ( n12 ) , .Y ( n10 ) ) ;
OAI21X1 U14 (.A ( alu_op[1] ) , .B ( alu_op[0] ) , .C ( n10 ) , .Y ( op[5] ) ) ;
NAND2X1 U13 (.A ( funct[1] ) , .B ( funct[0] ) , .Y ( n8 ) ) ;
NAND2X1 U12 (.A ( funct[2] ) , .B ( n4 ) , .Y ( n9 ) ) ;
OAI21X1 U11 (.A ( n8 ) , .B ( n9 ) , .C ( n1 ) , .Y ( op[6] ) ) ;
OR2X1 U26 (.A ( funct[0] ) , .B ( funct[2] ) , .Y ( n20 ) ) ;
NAND2X1 U25 (.A ( n4 ) , .B ( funct[1] ) , .Y ( n21 ) ) ;
AOI21X1 U24 (.A ( n2 ) , .B ( alu_op[0] ) , .C ( op[1] ) , .Y ( n16 ) ) ;
OAI21X1 U23 (.A ( n20 ) , .B ( n21 ) , .C ( n16 ) , .Y ( op[2] ) ) ;
NAND3X1 U22 (.A ( n19 ) , .B ( n7 ) , .C ( n11 ) , .Y ( n18 ) ) ;
OAI21X1 U21 (.A ( alu_op[1] ) , .B ( alu_op[0] ) , .C ( n18 ) , .Y ( op[3] ) ) ;
NAND3X1 U20 (.A ( funct[0] ) , .B ( n7 ) , .C ( funct[2] ) , .Y ( n14 ) ) ;
OAI21X1 U19 (.A ( n7 ) , .B ( funct[0] ) , .C ( n14 ) , .Y ( n17 ) ) ;
NOR2X1 U34 (.A ( funct[4] ) , .B ( alu_op[0] ) , .Y ( n26 ) ) ;
NAND2X1 U33 (.A ( n26 ) , .B ( funct[5] ) , .Y ( n25 ) ) ;
NOR2X1 U32 (.A ( n25 ) , .B ( funct[3] ) , .Y ( n11 ) ) ;
NAND2X1 U31 (.A ( n11 ) , .B ( alu_op[1] ) , .Y ( n15 ) ) ;
NAND2X1 U30 (.A ( funct[0] ) , .B ( n6 ) , .Y ( n19 ) ) ;
NOR2X1 U29 (.A ( n19 ) , .B ( n25 ) , .Y ( n23 ) ) ;
NAND3X1 U28 (.A ( n23 ) , .B ( alu_op[1] ) , .C ( n24 ) , .Y ( n22 ) ) ;
OAI21X1 U27 (.A ( n15 ) , .B ( n6 ) , .C ( n22 ) , .Y ( op[0] ) ) ;
endmodule


                                                                                                                                                                                                                       alu_ctl.pnr.v                                                                                       0000644 �    Asz0000145 00000013511 13055352430 011405  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   //
// Milkyway Hierarchical Verilog Dump:
// Generated on 02/28/2017 at 14:52:56
// Design Generated by Consolidated Verilog Reader
// File produced by Consolidated Verilog Writer
// Library Name :alu_ctl_LIB
// Cell Name    :alu_ctl
// Hierarchy delimiter:'/'
// Write Command : write_verilog alu_ctl.pnr.v
//


module alu_ctl (funct , alu_op , op );
input  [5:0] funct ;
input  [1:0] alu_op ;
output [6:0] op ;



INVX2 U10 (.A ( funct[1] ) , .Y ( n7 ) ) ;
INVX2 U9 (.A ( funct[2] ) , .Y ( n6 ) ) ;
INVX2 U8 (.A ( n17 ) , .Y ( n5 ) ) ;
INVX2 U7 (.A ( n15 ) , .Y ( n4 ) ) ;
INVX2 U6 (.A ( n22 ) , .Y ( op[1] ) ) ;
INVX2 U5 (.A ( alu_op[1] ) , .Y ( n2 ) ) ;
INVX2 U4 (.A ( op[2] ) , .Y ( n1 ) ) ;
AND2X2 U3 (.A ( funct[1] ) , .B ( funct[3] ) , .Y ( n24 ) ) ;
OAI21X1 U18 (.A ( n5 ) , .B ( n15 ) , .C ( n16 ) , .Y ( op[4] ) ) ;
XOR2X1 U17 (.A ( funct[2] ) , .B ( funct[1] ) , .Y ( n13 ) ) ;
OAI21X1 U16 (.A ( funct[0] ) , .B ( n13 ) , .C ( n14 ) , .Y ( n12 ) ) ;
NAND2X1 U15 (.A ( n11 ) , .B ( n12 ) , .Y ( n10 ) ) ;
OAI21X1 U14 (.A ( alu_op[1] ) , .B ( alu_op[0] ) , .C ( n10 ) , .Y ( op[5] ) ) ;
NAND2X1 U13 (.A ( funct[1] ) , .B ( funct[0] ) , .Y ( n8 ) ) ;
NAND2X1 U12 (.A ( funct[2] ) , .B ( n4 ) , .Y ( n9 ) ) ;
OAI21X1 U11 (.A ( n8 ) , .B ( n9 ) , .C ( n1 ) , .Y ( op[6] ) ) ;
OR2X1 U26 (.A ( funct[0] ) , .B ( funct[2] ) , .Y ( n20 ) ) ;
NAND2X1 U25 (.A ( n4 ) , .B ( funct[1] ) , .Y ( n21 ) ) ;
AOI21X1 U24 (.A ( n2 ) , .B ( alu_op[0] ) , .C ( op[1] ) , .Y ( n16 ) ) ;
OAI21X1 U23 (.A ( n20 ) , .B ( n21 ) , .C ( n16 ) , .Y ( op[2] ) ) ;
NAND3X1 U22 (.A ( n19 ) , .B ( n7 ) , .C ( n11 ) , .Y ( n18 ) ) ;
OAI21X1 U21 (.A ( alu_op[1] ) , .B ( alu_op[0] ) , .C ( n18 ) , .Y ( op[3] ) ) ;
NAND3X1 U20 (.A ( funct[0] ) , .B ( n7 ) , .C ( funct[2] ) , .Y ( n14 ) ) ;
OAI21X1 U19 (.A ( n7 ) , .B ( funct[0] ) , .C ( n14 ) , .Y ( n17 ) ) ;
NOR2X1 U34 (.A ( funct[4] ) , .B ( alu_op[0] ) , .Y ( n26 ) ) ;
NAND2X1 U33 (.A ( n26 ) , .B ( funct[5] ) , .Y ( n25 ) ) ;
NOR2X1 U32 (.A ( n25 ) , .B ( funct[3] ) , .Y ( n11 ) ) ;
NAND2X1 U31 (.A ( n11 ) , .B ( alu_op[1] ) , .Y ( n15 ) ) ;
NAND2X1 U30 (.A ( funct[0] ) , .B ( n6 ) , .Y ( n19 ) ) ;
NOR2X1 U29 (.A ( n19 ) , .B ( n25 ) , .Y ( n23 ) ) ;
NAND3X1 U28 (.A ( n23 ) , .B ( alu_op[1] ) , .C ( n24 ) , .Y ( n22 ) ) ;
OAI21X1 U27 (.A ( n15 ) , .B ( n6 ) , .C ( n22 ) , .Y ( op[0] ) ) ;
FILL xofiller_FILL_1 () ;
FILL xofiller_FILL_2 () ;
FILL xofiller_FILL_3 () ;
FILL xofiller_FILL_4 () ;
FILL xofiller_FILL_5 () ;
FILL xofiller_FILL_6 () ;
FILL xofiller_FILL_7 () ;
FILL xofiller_FILL_8 () ;
FILL xofiller_FILL_9 () ;
FILL xofiller_FILL_10 () ;
FILL xofiller_FILL_11 () ;
FILL xofiller_FILL_12 () ;
FILL xofiller_FILL_13 () ;
FILL xofiller_FILL_14 () ;
FILL xofiller_FILL_15 () ;
FILL xofiller_FILL_16 () ;
FILL xofiller_FILL_17 () ;
FILL xofiller_FILL_18 () ;
FILL xofiller_FILL_19 () ;
FILL xofiller_FILL_20 () ;
FILL xofiller_FILL_21 () ;
FILL xofiller_FILL_22 () ;
FILL xofiller_FILL_23 () ;
FILL xofiller_FILL_24 () ;
FILL xofiller_FILL_25 () ;
FILL xofiller_FILL_26 () ;
FILL xofiller_FILL_27 () ;
FILL xofiller_FILL_28 () ;
FILL xofiller_FILL_29 () ;
FILL xofiller_FILL_30 () ;
FILL xofiller_FILL_31 () ;
FILL xofiller_FILL_32 () ;
FILL xofiller_FILL_33 () ;
FILL xofiller_FILL_34 () ;
FILL xofiller_FILL_35 () ;
FILL xofiller_FILL_36 () ;
FILL xofiller_FILL_37 () ;
FILL xofiller_FILL_38 () ;
FILL xofiller_FILL_39 () ;
FILL xofiller_FILL_40 () ;
FILL xofiller_FILL_41 () ;
FILL xofiller_FILL_42 () ;
FILL xofiller_FILL_43 () ;
FILL xofiller_FILL_44 () ;
FILL xofiller_FILL_45 () ;
FILL xofiller_FILL_46 () ;
FILL xofiller_FILL_47 () ;
FILL xofiller_FILL_48 () ;
FILL xofiller_FILL_49 () ;
FILL xofiller_FILL_50 () ;
FILL xofiller_FILL_51 () ;
FILL xofiller_FILL_52 () ;
FILL xofiller_FILL_53 () ;
FILL xofiller_FILL_54 () ;
FILL xofiller_FILL_55 () ;
FILL xofiller_FILL_56 () ;
FILL xofiller_FILL_57 () ;
FILL xofiller_FILL_58 () ;
FILL xofiller_FILL_59 () ;
FILL xofiller_FILL_60 () ;
FILL xofiller_FILL_61 () ;
FILL xofiller_FILL_62 () ;
FILL xofiller_FILL_63 () ;
FILL xofiller_FILL_64 () ;
FILL xofiller_FILL_65 () ;
FILL xofiller_FILL_66 () ;
FILL xofiller_FILL_67 () ;
FILL xofiller_FILL_68 () ;
FILL xofiller_FILL_69 () ;
FILL xofiller_FILL_70 () ;
FILL xofiller_FILL_71 () ;
FILL xofiller_FILL_72 () ;
FILL xofiller_FILL_73 () ;
FILL xofiller_FILL_74 () ;
FILL xofiller_FILL_75 () ;
FILL xofiller_FILL_76 () ;
FILL xofiller_FILL_77 () ;
FILL xofiller_FILL_78 () ;
FILL xofiller_FILL_79 () ;
FILL xofiller_FILL_80 () ;
FILL xofiller_FILL_81 () ;
FILL xofiller_FILL_82 () ;
FILL xofiller_FILL_83 () ;
FILL xofiller_FILL_84 () ;
FILL xofiller_FILL_85 () ;
FILL xofiller_FILL_86 () ;
FILL xofiller_FILL_87 () ;
FILL xofiller_FILL_88 () ;
FILL xofiller_FILL_89 () ;
FILL xofiller_FILL_90 () ;
FILL xofiller_FILL_91 () ;
FILL xofiller_FILL_92 () ;
FILL xofiller_FILL_93 () ;
FILL xofiller_FILL_94 () ;
FILL xofiller_FILL_95 () ;
FILL xofiller_FILL_96 () ;
FILL xofiller_FILL_97 () ;
FILL xofiller_FILL_98 () ;
FILL xofiller_FILL_99 () ;
FILL xofiller_FILL_100 () ;
FILL xofiller_FILL_101 () ;
FILL xofiller_FILL_102 () ;
FILL xofiller_FILL_103 () ;
FILL xofiller_FILL_104 () ;
FILL xofiller_FILL_105 () ;
FILL xofiller_FILL_106 () ;
FILL xofiller_FILL_107 () ;
FILL xofiller_FILL_108 () ;
FILL xofiller_FILL_109 () ;
FILL xofiller_FILL_110 () ;
FILL xofiller_FILL_111 () ;
FILL xofiller_FILL_112 () ;
FILL xofiller_FILL_113 () ;
FILL xofiller_FILL_114 () ;
FILL xofiller_FILL_115 () ;
FILL xofiller_FILL_116 () ;
FILL xofiller_FILL_117 () ;
FILL xofiller_FILL_118 () ;
FILL xofiller_FILL_119 () ;
FILL xofiller_FILL_120 () ;
FILL xofiller_FILL_121 () ;
FILL xofiller_FILL_122 () ;
FILL xofiller_FILL_123 () ;
FILL xofiller_FILL_124 () ;
FILL xofiller_FILL_125 () ;
FILL xofiller_FILL_126 () ;
FILL xofiller_FILL_127 () ;
FILL xofiller_FILL_128 () ;
FILL xofiller_FILL_129 () ;
FILL xofiller_FILL_130 () ;
FILL xofiller_FILL_131 () ;
FILL xofiller_FILL_132 () ;
FILL xofiller_FILL_133 () ;
endmodule


                                                                                                                                                                                       alu_ctl.post_synth.v                                                                                0000644 �    Asz0000145 00000004075 13055347052 013031  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   /////////////////////////////////////////////////////////////
// Created by: Synopsys DC Expert(TM) in wire load mode
// Version   : L-2016.03-SP5-2
// Date      : Tue Feb 28 14:23:22 2017
/////////////////////////////////////////////////////////////


module alu_ctl ( alu_op, funct, op );
  input [1:0] alu_op;
  input [5:0] funct;
  output [6:0] op;
  wire   n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  AND2X2 U3 ( .A(funct[1]), .B(funct[3]), .Y(n24) );
  INVX2 U4 ( .A(op[2]), .Y(n1) );
  INVX2 U5 ( .A(alu_op[1]), .Y(n2) );
  INVX2 U6 ( .A(n22), .Y(op[1]) );
  INVX2 U7 ( .A(n15), .Y(n4) );
  INVX2 U8 ( .A(n17), .Y(n5) );
  INVX2 U9 ( .A(funct[2]), .Y(n6) );
  INVX2 U10 ( .A(funct[1]), .Y(n7) );
  OAI21X1 U11 ( .A(n8), .B(n9), .C(n1), .Y(op[6]) );
  NAND2X1 U12 ( .A(funct[2]), .B(n4), .Y(n9) );
  NAND2X1 U13 ( .A(funct[1]), .B(funct[0]), .Y(n8) );
  OAI21X1 U14 ( .A(alu_op[1]), .B(alu_op[0]), .C(n10), .Y(op[5]) );
  NAND2X1 U15 ( .A(n11), .B(n12), .Y(n10) );
  OAI21X1 U16 ( .A(funct[0]), .B(n13), .C(n14), .Y(n12) );
  XOR2X1 U17 ( .A(funct[2]), .B(funct[1]), .Y(n13) );
  OAI21X1 U18 ( .A(n5), .B(n15), .C(n16), .Y(op[4]) );
  OAI21X1 U19 ( .A(n7), .B(funct[0]), .C(n14), .Y(n17) );
  NAND3X1 U20 ( .A(funct[0]), .B(n7), .C(funct[2]), .Y(n14) );
  OAI21X1 U21 ( .A(alu_op[1]), .B(alu_op[0]), .C(n18), .Y(op[3]) );
  NAND3X1 U22 ( .A(n19), .B(n7), .C(n11), .Y(n18) );
  OAI21X1 U23 ( .A(n20), .B(n21), .C(n16), .Y(op[2]) );
  AOI21X1 U24 ( .A(n2), .B(alu_op[0]), .C(op[1]), .Y(n16) );
  NAND2X1 U25 ( .A(n4), .B(funct[1]), .Y(n21) );
  OR2X1 U26 ( .A(funct[0]), .B(funct[2]), .Y(n20) );
  OAI21X1 U27 ( .A(n15), .B(n6), .C(n22), .Y(op[0]) );
  NAND3X1 U28 ( .A(n23), .B(alu_op[1]), .C(n24), .Y(n22) );
  NOR2X1 U29 ( .A(n19), .B(n25), .Y(n23) );
  NAND2X1 U30 ( .A(funct[0]), .B(n6), .Y(n19) );
  NAND2X1 U31 ( .A(n11), .B(alu_op[1]), .Y(n15) );
  NOR2X1 U32 ( .A(n25), .B(funct[3]), .Y(n11) );
  NAND2X1 U33 ( .A(n26), .B(funct[5]), .Y(n25) );
  NOR2X1 U34 ( .A(funct[4]), .B(alu_op[0]), .Y(n26) );
endmodule

                                                                                                                                                                                                                                                                                                                                                                                                                                                                   counter_bench.v                                                                                     0000644 �    Asz0000145 00000001313 12317616736 012013  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   module counter_bench;
   reg clk, clr, up;
   wire [3:0] Q;
   
   counter DUV (clk, clr, up, Q);

   always begin
      clk = 0;
      #10;
      clk = 1;
      #10;
   end

   initial begin
      $vcdpluson;   /* dump signals to file vcdplus.vcd */
      clr = 1;
      up = 0;
      #1;
      @(posedge clk) #1;
      clr = 0;
      $display("time=%t, clr=%d, up=%d, Q=%h", $time, clr, up, Q);
      repeat (18) begin
	 @(posedge clk) #1;
	 $display("time=%t, clr=%d, up=%d, Q=%h", $time, clr, up, Q);
      end
      up = 1;
      repeat (18) begin
	 @(posedge clk) #1;
	 $display("time=%t, clr=%d, up=%d, Q=%h", $time, clr, up, Q);
      end
      $finish;
   end // initial begin
endmodule // counter_bench


                                                                                                                                                                                                                                                                                                                     counter.v                                                                                           0000644 �    Asz0000145 00000000532 12317072532 010644  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   module counter(input clk, input clr, input up,
	       output reg [3:0] Q /*, output carry*/);



//   assign 	      carry =  ( up && (Q == 4'b1111) )
//                            || (~up && (Q == 4'b0000));
   
   always @(posedge clk)
     begin
	if (clr) Q <= 4'd0;
	else if (up) Q <= Q + 1;
	else Q <= Q - 1;
     end

endmodule // counter

                                                                                                                                                                      decoder_bench.v                                                                                     0000644 �    Asz0000145 00000001436 12317355312 011735  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   module decoder_bench;

   reg [1:0] a;
   wire      y0, y1, y2, y3;
   
   decoder DUV (a, y0, y1, y2, y3);

   initial begin
      $vcdpluson;   /* dump signals to file vcdplus.vcd */
      a = 2'd0;
      #10;       
      $display("time=%t a=%d y0y1y2y3 = %b %b %b %b", $time, a, y0, y1, y2, y3);
      a = 2'd1;
      #10;
      $display("time=%t a=%d y0y1y2y3 = %b %b %b %b", $time, a, y0, y1, y2, y3);
      a = 2'd2;
      #10;
      $display("time=%t a=%d y0y1y2y3 = %b %b %b %b", $time, a, y0, y1, y2, y3);
      a = 2'd3;
      #10;
      $display("time=%t a=%d y0y1y2y3 = %b %b %b %b", $time, a, y0, y1, y2, y3);
      a = 2'd0;
      #10;
      $display("time=%t a=%d y0y1y2y3 = %b %b %b %b", $time, a, y0, y1, y2, y3);
      $finish;
   end // initial begin
endmodule // decoder_test

                                                                                                                                                                                                                                  decoder.nofill.v                                                                                    0000644 �    Asz0000145 00000001312 13055336335 012055  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   //
// Milkyway Hierarchical Verilog Dump:
// Generated on 02/28/2017 at 13:09:33
// Design Generated by Consolidated Verilog Reader
// File produced by Consolidated Verilog Writer
// Library Name :decoder_LIB
// Cell Name    :decoder
// Hierarchy delimiter:'/'
// Write Command : write_verilog decoder.pnr.v
//


module decoder (y3 , y2 , y1 , y0 , a );
output y3 ;
output y2 ;
output y1 ;
output y0 ;
input  [1:0] a ;



NOR2X1 U8 (.A ( a[1] ) , .B ( a[0] ) , .Y ( y0 ) ) ;
NOR2X1 U7 (.A ( a[1] ) , .B ( n2 ) , .Y ( y1 ) ) ;
NOR2X1 U6 (.A ( a[0] ) , .B ( n1 ) , .Y ( y2 ) ) ;
NOR2X1 U5 (.A ( n2 ) , .B ( n1 ) , .Y ( y3 ) ) ;
INVX2 U4 (.A ( a[0] ) , .Y ( n2 ) ) ;
INVX2 U3 (.A ( a[1] ) , .Y ( n1 ) ) ;
endmodule


                                                                                                                                                                                                                                                                                                                      decoder.pnr.v                                                                                       0000644 �    Asz0000145 00000002126 13055336335 011375  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   //
// Milkyway Hierarchical Verilog Dump:
// Generated on 02/28/2017 at 13:09:33
// Design Generated by Consolidated Verilog Reader
// File produced by Consolidated Verilog Writer
// Library Name :decoder_LIB
// Cell Name    :decoder
// Hierarchy delimiter:'/'
// Write Command : write_verilog decoder.pnr.v
//


module decoder (y3 , y2 , y1 , y0 , a );
output y3 ;
output y2 ;
output y1 ;
output y0 ;
input  [1:0] a ;



NOR2X1 U8 (.A ( a[1] ) , .B ( a[0] ) , .Y ( y0 ) ) ;
NOR2X1 U7 (.A ( a[1] ) , .B ( n2 ) , .Y ( y1 ) ) ;
NOR2X1 U6 (.A ( a[0] ) , .B ( n1 ) , .Y ( y2 ) ) ;
NOR2X1 U5 (.A ( n2 ) , .B ( n1 ) , .Y ( y3 ) ) ;
INVX2 U4 (.A ( a[0] ) , .Y ( n2 ) ) ;
INVX2 U3 (.A ( a[1] ) , .Y ( n1 ) ) ;
FILL xofiller_FILL_1 () ;
FILL xofiller_FILL_2 () ;
FILL xofiller_FILL_3 () ;
FILL xofiller_FILL_4 () ;
FILL xofiller_FILL_5 () ;
FILL xofiller_FILL_6 () ;
FILL xofiller_FILL_7 () ;
FILL xofiller_FILL_8 () ;
FILL xofiller_FILL_9 () ;
FILL xofiller_FILL_10 () ;
FILL xofiller_FILL_11 () ;
FILL xofiller_FILL_12 () ;
FILL xofiller_FILL_13 () ;
FILL xofiller_FILL_14 () ;
FILL xofiller_FILL_15 () ;
endmodule


                                                                                                                                                                                                                                                                                                                                                                                                                                          decoder.post_synth.v                                                                                0000644 �    Asz0000145 00000001124 13055346456 013012  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   /////////////////////////////////////////////////////////////
// Created by: Synopsys DC Expert(TM) in wire load mode
// Version   : L-2016.03-SP5-2
// Date      : Tue Feb 28 14:19:10 2017
/////////////////////////////////////////////////////////////


module decoder ( a, y0, y1, y2, y3 );
  input [1:0] a;
  output y0, y1, y2, y3;
  wire   n1, n2;

  INVX2 U3 ( .A(a[1]), .Y(n1) );
  INVX2 U4 ( .A(a[0]), .Y(n2) );
  NOR2X1 U5 ( .A(n2), .B(n1), .Y(y3) );
  NOR2X1 U6 ( .A(a[0]), .B(n1), .Y(y2) );
  NOR2X1 U7 ( .A(a[1]), .B(n2), .Y(y1) );
  NOR2X1 U8 ( .A(a[1]), .B(a[0]), .Y(y0) );
endmodule

                                                                                                                                                                                                                                                                                                                                                                                                                                            decoder.v                                                                                           0000644 �    Asz0000145 00000000516 12317072436 010577  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   module decoder(a,y0,y1,y2,y3);
   input [1:0] a;
   output      y0, y1, y2, y3;
   reg 	       y0, y1, y2, y3;

   always @(a)
      begin
	 y0 = 0;
	 y1 = 0;
	 y2 = 0;
	 y3 = 0;
	 case (a)
	   2'b00: y0 = 1;
	   2'b01: y1 = 1;
	   2'b10: y2 = 1;
	   2'b11: y3 = 1;
	 endcase // case(a)
      end // always @ (a)
endmodule // decoder
                                                                                                                                                                                  iccscript_comb_new.tcl                                                                              0000644 �    Asz0000145 00000010400 13055352364 013335  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   ############################################################################
# ON C5 0.5u CMOS ASIC Place and Route Script using IC Compiler - Version 3.0
#############################################################################
# This script assumes that the post synthesis netlist and sdc file produced by 
#   synthesis are both in the local directory
#############################################################################
# Update the lib_path and design_name for your design
#############################################################################
set OSUcells "/home/shared/OSU/synopsys/lib/ami05"
#set OSUcells [format "%s%s"  [getenv "OSUcells"] "/lib/ami05"]
#set         lib_path    "/users/eesunz/faculty/cdsemac/UofU_SYNS_v1_2/UTFSM_libraries"
set         lib_path    $OSUcells

## modify design_name to match your design
set         design_name    "alu_ctl"  

set_app_var search_path "$lib_path"
set_app_var target_library "osu05_stdcells.db"
set_app_var link_library "* $target_library"

#if { ( file exists "[set design_name]_LIB" ) } { sh rm -rf "[set design_name]_LIB" }
sh rm -rf ${design_name}_LIB

create_mw_lib -tech "/home/shared/OSU/synopsys/flow/ami05/tech.tf" -mw_reference_library "$lib_path/osu05_stdcells"  ${design_name}_LIB

open_mw_lib   "${design_name}_LIB"

#set_tlu_plus_files  \
#    -max_tluplus  "$lib_path/MW_UTAH/ami500.tluplus"   \
#    -min_tluplus  "$lib_path/MW_UTAH/ami500.tluplus"   \
#    -tech2itf_map "$lib_path/MW_UTAH/ami500hxkx_3m.map"

import_design   "./${design_name}.post_synth.v"  -format "verilog" -top ${design_name} -cel ${design_name} 

read_sdc ./${design_name}.sdc

#### Add pin constraints here to set pin placement
#  Note that sides are numbered as follows:
#    side 1: LEFT
#    side 2: TOP
#    side 3: RIGHT
#    side 4: BOTTOM
#  the offset value is in microns starting from the lower coordinate of the referenced side
#
#  As an example, the following will place a pin named "myPin" on the bottom of the cell
#  10 microns from its left edge:
# set_pin_physical_constraints -pin_name {myPin} -layers {metal2} -side 4 -offset 10

###### Adjust density here to alleviate LVS errors after routing at the expense of a larger design
create_floorplan -control_type "aspect_ratio" -core_aspect_ratio "3.5" -core_utilization "0.4" -row_core_ratio "1" -start_first_row  -left_io2core 24 -bottom_io2core 27 -right_io2core 24 -top_io2core 27

derive_pg_connection -power_net {vdd!} -ground_net {gnd!}

create_rectilinear_rings -nets {vdd! gnd!} -offset {3 3} -width {4.5 4.5} -space {3 3}

###### Adjust the number of straps here to alleviate LVS problems after routing  - at the expense of a less robust power network
create_power_straps  -direction vertical -num_placement_strap 1 -start_at 400 -increment_x_or_y 200 -nets  {vdd! gnd!}  -width 1.800 -layer metal3

place_opt -effort high -congestion

preroute_standard_cells -nets {vdd! gnd!} -connect horizontal -extend_to_boundaries_and_generate_pins 

#clock_opt -fix_hold_all_clocks

#report_clock_tree

report_timing

route_zrt_auto -max_detail_route_iterations 1000
route_zrt_detail -incremental true

insert_stdcell_filler -cell_without_metal "FILL8 FILL4 FILL2 FILL"  -connect_to_power "vdd!" -connect_to_ground "gnd!"

preroute_standard_cells -nets {vdd! gnd!} -connect horizontal -extend_to_boundaries_and_generate_pins 

derive_pg_connection -power_net {vdd!} -ground_net {gnd!}

# This command shows a warning that the command is old and no longer valid.
# Not really true.  For designs in deep submicron (65nm and below) you should use the new checker.
# However for designs older than 65nm, this is the appropriate checker.   

verify_drc

verify_lvs

route_zrt_detail -incremental true

report_timing > ${design_name}.timing

change_names -rules verilog -hierarchy

write_verilog ${design_name}.pnr.v

sh grep -v FILL ${design_name}.pnr.v > ${design_name}.nofill.v 


set_write_stream_options -output_pin {text geometry} -keep_data_type -child_depth 20 -map_layer "/home/shared/OSU/synopsys/flow/ami05/streamout.map"
write_stream -lib_name ${design_name}_LIB -format gds ${design_name}.gds

write_sdc     ${design_name}.pnr.sdc

extract_rc -coupling_cap

write_parasitics -format SBPF -output "${design_name}.pnr.sbpf"

verify_pg_nets

report_timing 

#report_clock_tree

save_mw_cel

##close_mw_cel

##exit
                                                                                                                                                                                                                                                                iccscript_comb_orig.tcl                                                                             0000644 �    Asz0000145 00000007360 13051117406 013507  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   ############################################################################
# ON C5 0.5u CMOS ASIC Place and Route Script using IC Compiler - Version 3.0
#############################################################################
# This script assumes that the post synthesis netlist and sdc file produced by 
#   synthesis are both in the local directory
#############################################################################
# Update the lib_path and design_name for your design
#############################################################################
set OSUcells [format "%s%s"  [getenv "OSUcells"] "/lib/ami05"]
#set         lib_path    "/users/eesunz/faculty/cdsemac/UofU_SYNS_v1_2/UTFSM_libraries"
set         lib_path    $OSUcells

## modify design_name to match your design
set         design_name    "decoder"  

set_app_var search_path "$lib_path"
set_app_var target_library "osu05_stdcells.db"
set_app_var link_library "* $target_library"

#if { ( file exists "[set design_name]_LIB" ) } { sh rm -rf "[set design_name]_LIB" }
sh rm -rf ${design_name}_LIB

create_mw_lib -tech "/usr14/cad/OSU/synopsys/flow/ami05/tech.tf" -mw_reference_library "$lib_path/osu05_stdcells"  ${design_name}_LIB

open_mw_lib   "${design_name}_LIB"

#set_tlu_plus_files  \
#    -max_tluplus  "$lib_path/MW_UTAH/ami500.tluplus"   \
#    -min_tluplus  "$lib_path/MW_UTAH/ami500.tluplus"   \
#    -tech2itf_map "$lib_path/MW_UTAH/ami500hxkx_3m.map"

import_design   "./${design_name}.post_synth.v"  -format "verilog" -top ${design_name} -cel ${design_name} 

read_sdc ./${design_name}.sdc

###### Adjust density here to alleviate LVS errors after routing at the expense of a larger design
create_floorplan -control_type "aspect_ratio" -core_aspect_ratio "0.5" -core_utilization "0.4" -row_core_ratio "1" -start_first_row  -left_io2core 24 -bottom_io2core 27 -right_io2core 24 -top_io2core 27

derive_pg_connection -power_net {vdd!} -ground_net {gnd!}

create_rectilinear_rings -nets {vdd! gnd!} -offset {3 3} -width {4.5 4.5} -space {3 3}

###### Adjust the number of straps here to alleviate LVS problems after routing  - at the expense of a less robust power network
create_power_straps  -direction vertical -num_placement_strap 1 -start_at 400 -increment_x_or_y 200 -nets  {vdd! gnd!}  -width 1.800 -layer metal3

place_opt -effort high -congestion

preroute_standard_cells -nets {vdd! gnd!} -connect horizontal -extend_to_boundaries_and_generate_pins 

#clock_opt -fix_hold_all_clocks

#report_clock_tree

report_timing

route_zrt_auto -max_detail_route_iterations 1000
route_zrt_detail -incremental true

insert_stdcell_filler -cell_without_metal "FILL8 FILL4 FILL2 FILL"  -connect_to_power "vdd!" -connect_to_ground "gnd!"

preroute_standard_cells -nets {vdd! gnd!} -connect horizontal -extend_to_boundaries_and_generate_pins 

derive_pg_connection -power_net {vdd!} -ground_net {gnd!}

# This command shows a warning that the command is old and no longer valid.
# Not really true.  For designs in deep submicron (65nm and below) you should use the new checker.
# However for designs older than 65nm, this is the appropriate checker.   

verify_drc

verify_lvs

route_zrt_detail -incremental true

report_timing > ${design_name}.timing

change_names -rules verilog -hierarchy

write_verilog ${design_name}.pnr.v

sh grep -v FILL ${design_name}.pnr.v > ${design_name}.nofill.v 


set_write_stream_options -output_pin {text geometry} -keep_data_type -child_depth 20 -map_layer "/usr14/cad/OSU/synopsys/flow/ami05/streamout.map"
write_stream -lib_name ${design_name}_LIB -format gds ${design_name}.gds

write_sdc     ${design_name}.pnr.sdc

extract_rc -coupling_cap

write_parasitics -format SBPF -output "${design_name}.pnr.sbpf"

verify_pg_nets

report_timing 

#report_clock_tree

save_mw_cel

##close_mw_cel

##exit
                                                                                                                                                                                                                                                                                iccscript_comb.tcl                                                                                  0000644 �    Asz0000145 00000010400 13054651325 012462  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   ############################################################################
# ON C5 0.5u CMOS ASIC Place and Route Script using IC Compiler - Version 3.0
#############################################################################
# This script assumes that the post synthesis netlist and sdc file produced by 
#   synthesis are both in the local directory
#############################################################################
# Update the lib_path and design_name for your design
#############################################################################
set OSUcells "/home/shared/OSU/synopsys/lib/ami05"
#set OSUcells [format "%s%s"  [getenv "OSUcells"] "/lib/ami05"]
#set         lib_path    "/users/eesunz/faculty/cdsemac/UofU_SYNS_v1_2/UTFSM_libraries"
set         lib_path    $OSUcells

## modify design_name to match your design
set         design_name    "decoder"  

set_app_var search_path "$lib_path"
set_app_var target_library "osu05_stdcells.db"
set_app_var link_library "* $target_library"

#if { ( file exists "[set design_name]_LIB" ) } { sh rm -rf "[set design_name]_LIB" }
sh rm -rf ${design_name}_LIB

create_mw_lib -tech "/home/shared/OSU/synopsys/flow/ami05/tech.tf" -mw_reference_library "$lib_path/osu05_stdcells"  ${design_name}_LIB

open_mw_lib   "${design_name}_LIB"

#set_tlu_plus_files  \
#    -max_tluplus  "$lib_path/MW_UTAH/ami500.tluplus"   \
#    -min_tluplus  "$lib_path/MW_UTAH/ami500.tluplus"   \
#    -tech2itf_map "$lib_path/MW_UTAH/ami500hxkx_3m.map"

import_design   "./${design_name}.post_synth.v"  -format "verilog" -top ${design_name} -cel ${design_name} 

read_sdc ./${design_name}.sdc

#### Add pin constraints here to set pin placement
#  Note that sides are numbered as follows:
#    side 1: LEFT
#    side 2: TOP
#    side 3: RIGHT
#    side 4: BOTTOM
#  the offset value is in microns starting from the lower coordinate of the referenced side
#
#  As an example, the following will place a pin named "myPin" on the bottom of the cell
#  10 microns from its left edge:
# set_pin_physical_constraints -pin_name {myPin} -layers {metal2} -side 4 -offset 10

###### Adjust density here to alleviate LVS errors after routing at the expense of a larger design
create_floorplan -control_type "aspect_ratio" -core_aspect_ratio "0.5" -core_utilization "0.4" -row_core_ratio "1" -start_first_row  -left_io2core 24 -bottom_io2core 27 -right_io2core 24 -top_io2core 27

derive_pg_connection -power_net {vdd!} -ground_net {gnd!}

create_rectilinear_rings -nets {vdd! gnd!} -offset {3 3} -width {4.5 4.5} -space {3 3}

###### Adjust the number of straps here to alleviate LVS problems after routing  - at the expense of a less robust power network
create_power_straps  -direction vertical -num_placement_strap 1 -start_at 400 -increment_x_or_y 200 -nets  {vdd! gnd!}  -width 1.800 -layer metal3

place_opt -effort high -congestion

preroute_standard_cells -nets {vdd! gnd!} -connect horizontal -extend_to_boundaries_and_generate_pins 

#clock_opt -fix_hold_all_clocks

#report_clock_tree

report_timing

route_zrt_auto -max_detail_route_iterations 1000
route_zrt_detail -incremental true

insert_stdcell_filler -cell_without_metal "FILL8 FILL4 FILL2 FILL"  -connect_to_power "vdd!" -connect_to_ground "gnd!"

preroute_standard_cells -nets {vdd! gnd!} -connect horizontal -extend_to_boundaries_and_generate_pins 

derive_pg_connection -power_net {vdd!} -ground_net {gnd!}

# This command shows a warning that the command is old and no longer valid.
# Not really true.  For designs in deep submicron (65nm and below) you should use the new checker.
# However for designs older than 65nm, this is the appropriate checker.   

verify_drc

verify_lvs

route_zrt_detail -incremental true

report_timing > ${design_name}.timing

change_names -rules verilog -hierarchy

write_verilog ${design_name}.pnr.v

sh grep -v FILL ${design_name}.pnr.v > ${design_name}.nofill.v 


set_write_stream_options -output_pin {text geometry} -keep_data_type -child_depth 20 -map_layer "/home/shared/OSU/synopsys/flow/ami05/streamout.map"
write_stream -lib_name ${design_name}_LIB -format gds ${design_name}.gds

write_sdc     ${design_name}.pnr.sdc

extract_rc -coupling_cap

write_parasitics -format SBPF -output "${design_name}.pnr.sbpf"

verify_pg_nets

report_timing 

#report_clock_tree

save_mw_cel

##close_mw_cel

##exit
                                                                                                                                                                                                                                                                iccscript.tcl                                                                                       0000644 �    Asz0000145 00000010406 13054651321 011464  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   #############################################################################
# ON C5 0.5u CMOS ASIC Place and Route Script using IC Compiler - Version 3.0
#############################################################################
# This script assumes that the post synthesis netlist and sdc file produced by 
#   synthesis are both in the local directory
#############################################################################
# Update the lib_path and design_name for your design
#############################################################################
set OSUcells "/home/shared/OSU/synopsys/lib/ami05"
#set OSUcells [format "%s%s"  [getenv "OSUcells"] "synopsys/lib/ami05"]
#set         lib_path    "/users/eesunz/faculty/cdsemac/UofU_SYNS_v1_2/UTFSM_libraries"
set          lib_path    $OSUcells

## modify design_name to match your design
set         design_name    "counter"  

set_app_var search_path "$lib_path"
set_app_var target_library "osu05_stdcells.db"
set_app_var link_library "* $target_library"

#if { ( file exists "[set design_name]_LIB" ) } { sh rm -rf "[set design_name]_LIB" }
sh rm -rf ${design_name}_LIB

create_mw_lib -tech "/home/shared/OSU/synopsys/flow/ami05/tech.tf" -mw_reference_library "$lib_path/osu05_stdcells"  ${design_name}_LIB

open_mw_lib   "${design_name}_LIB"

#set_tlu_plus_files  \
#    -max_tluplus  "$lib_path/MW_UTAH/ami500.tluplus"   \
#    -min_tluplus  "$lib_path/MW_UTAH/ami500.tluplus"   \
#    -tech2itf_map "$lib_path/MW_UTAH/ami500hxkx_3m.map"

import_design   "./${design_name}.post_synth.v"  -format "verilog" -top ${design_name} -cel ${design_name} 

read_sdc ./${design_name}.sdc

#### Add pin constraints here to set pin placement
#  Note that sides are numbered as follows:
#    side 1: LEFT
#    side 2: TOP
#    side 3: RIGHT
#    side 4: BOTTOM
#  the offset value is in microns starting from the lower coordinate of the referenced side
#
#  As an example, the following will place a pin named "myPin" on the bottom of the cell
#  10 microns from its left edge:
# set_pin_physical_constraints -pin_name {myPin} -layers {metal2} -side 4 -offset 10

###### Adjust density here to alleviate LVS errors after routing at the expense of a larger design
create_floorplan -control_type "aspect_ratio" -core_aspect_ratio "0.5" -core_utilization "0.6" -row_core_ratio "1" -start_first_row  -left_io2core 24 -bottom_io2core 27 -right_io2core 24 -top_io2core 27

derive_pg_connection -power_net {vdd!} -ground_net {gnd!}

create_rectilinear_rings -nets {vdd! gnd!} -offset {3 3} -width {4.5 4.5} -space {3 3}

###### Adjust the number of straps here to alleviate LVS problems after routing  - at the expense of a less robust power network
create_power_straps  -direction vertical -num_placement_strap 1 -start_at 400 -increment_x_or_y 200 -nets  {vdd! gnd!}  -width 1.800 -layer metal3

place_opt -effort high -congestion

preroute_standard_cells -nets {vdd! gnd!} -connect horizontal -extend_to_boundaries_and_generate_pins 

clock_opt -fix_hold_all_clocks

report_clock_tree

report_timing

route_zrt_auto -max_detail_route_iterations 1000
route_zrt_detail -incremental true

insert_stdcell_filler -cell_without_metal "FILL8 FILL4 FILL2 FILL"  -connect_to_power "vdd!" -connect_to_ground "gnd!"

preroute_standard_cells -nets {vdd! gnd!} -connect horizontal -extend_to_boundaries_and_generate_pins 

derive_pg_connection -power_net {vdd!} -ground_net {gnd!}

# This command shows a warning that the command is old and no longer valid.
# Not really true.  For designs in deep submicron (65nm and below) you should use the new checker.
# However for designs older than 65nm, this is the appropriate checker.   

verify_drc

verify_lvs

route_zrt_detail -incremental true

report_timing > ${design_name}.timing

change_names -rules verilog -hierarchy

write_verilog ${design_name}.pnr.v

sh grep -v FILL ${design_name}.pnr.v > ${design_name}.nofill.v 

set_write_stream_options -output_pin {text geometry} -keep_data_type -child_depth 20 -map_layer "/home/shared/OSU/synopsys/flow/ami05/streamout.map"
write_stream -lib_name ${design_name}_LIB -format gds ${design_name}.gds

write_sdc     ${design_name}.pnr.sdc

extract_rc -coupling_cap

write_parasitics -format SBPF -output "${design_name}.pnr.sbpf"

verify_pg_nets

report_timing 

report_clock_tree

save_mw_cel

##close_mw_cel

##exit
                                                                                                                                                                                                                                                          synthesis_comb_new.tcl                                                                              0000644 �    Asz0000145 00000004741 13055347045 013416  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   #############################
# Script to synthesize combinational logic
# (customized from general script)
#############################

#############################
#  Change the following to your top-level design name
#############################

set         design_name    "alu_ctl"  

## hacked to work with OSU ami05 library - JN 3/27/14

set OSUcells "/home/shared/OSU/synopsys/lib/ami05"

set search_path [concat  $search_path $OSUcells]

set target_library [list osu05_stdcells.db]

set synthetic_library [list dw_foundation.sldb standard.sldb]

set link_library [concat $target_library $synthetic_library]

### following line stolen from OSU flow:
set alib_library_analysis_path $OSUcells

define_design_lib work -path ./work


#############################
# Read the verilog file.  If you use submodules,
# add commands to read thim first.
#############################
analyze -format sverilog ./${design_name}.sv

#############################
#  Translate the design into generic hardware
#############################
elaborate ${design_name}

#############################
# Set up clock and timing constratins
# Note that since there are no clocks in comb. logic
# clock constraints are commented out
#############################
set_max_delay 25 -to [all_outputs]
#create_clock "clk" -period 200
#create_clock "clk_in2" -period 100
#create_clock "clk_in3" -period 100

#############################
# if you have an internally generated clock instantiate a buffer (BUFX2)
# to provide a pin to identify the source of your new clock
#############################
#create_generated_clock -divide_by 1024 -source clk_in1 [get_pins {buffer/Y}]

#report_clocks

check_design > check_design.output

############################
# Make unique copies of submodules;
# Optimize & map to hardware
###########################
ungroup -flatten -all

set_flatten true -effort high
uniquify

compile

#############################
# Check these files once completed 
#############################
report_area  > area.rpt
report_hierarchy > hierarchy.rpt
report_constraints > constraints.rpt
report_timing > timing.rpt

#set_propagated_clock [all_clocks]

#############################
# Your timing file for IC Compiler 
#############################
write_sdc  ${design_name}.sdc

#############################
# Your output netlist 
#############################
write -f verilog ${design_name} -output ${design_name}.post_synth.v -hierarchy

# remove the comment if you want to leave dc_shell upon completion
# exit
                               synthesis_comb.tcl                                                                                  0000644 �    Asz0000145 00000004737 13051121350 012533  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   #############################
# Script to synthesize combinational logic
# (customized from general script)
#############################

#############################
#  Change the following to your top-level design name
#############################

set         design_name    "decoder"  

## hacked to work with OSU ami05 library - JN 3/27/14

set OSUcells "/home/shared/OSU/synopsys/lib/ami05"

set search_path [concat  $search_path $OSUcells]

set target_library [list osu05_stdcells.db]

set synthetic_library [list dw_foundation.sldb standard.sldb]

set link_library [concat $target_library $synthetic_library]

### following line stolen from OSU flow:
set alib_library_analysis_path $OSUcells

define_design_lib work -path ./work


#############################
# Read the verilog file.  If you use submodules,
# add commands to read thim first.
#############################
analyze -format verilog ./${design_name}.v

#############################
#  Translate the design into generic hardware
#############################
elaborate ${design_name}

#############################
# Set up clock and timing constratins
# Note that since there are no clocks in comb. logic
# clock constraints are commented out
#############################
set_max_delay 25 -to [all_outputs]
#create_clock "clk" -period 200
#create_clock "clk_in2" -period 100
#create_clock "clk_in3" -period 100

#############################
# if you have an internally generated clock instantiate a buffer (BUFX2)
# to provide a pin to identify the source of your new clock
#############################
#create_generated_clock -divide_by 1024 -source clk_in1 [get_pins {buffer/Y}]

#report_clocks

check_design > check_design.output

############################
# Make unique copies of submodules;
# Optimize & map to hardware
###########################
ungroup -flatten -all

set_flatten true -effort high
uniquify

compile

#############################
# Check these files once completed 
#############################
report_area  > area.rpt
report_hierarchy > hierarchy.rpt
report_constraints > constraints.rpt
report_timing > timing.rpt

#set_propagated_clock [all_clocks]

#############################
# Your timing file for IC Compiler 
#############################
write_sdc  ${design_name}.sdc

#############################
# Your output netlist 
#############################
write -f verilog ${design_name} -output ${design_name}.post_synth.v -hierarchy

# remove the comment if you want to leave dc_shell upon completion
# exit
                                 synthesis.tcl                                                                                       0000644 �    Asz0000145 00000004411 13053665170 011537  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   #############################
# Script to synthesize combinational logic
# (customized from general script)
#############################

#############################
#  Change the following to your top-level design name
#############################

set         design_name    "counter"  

## hacked to work with OSU ami05 library - JN 3/27/14

set OSUcells "/home/shared/OSU/synopsys/lib/ami05"

set search_path [concat  $search_path $OSUcells]

set target_library [list osu05_stdcells.db]

set synthetic_library [list dw_foundation.sldb standard.sldb]

set link_library [concat $target_library $synthetic_library]

### following line stolen from OSU flow:
set alib_library_analysis_path $OSUcells

define_design_lib work -path ./work


#############################
# Change this to your top-level file
# (include any other files containing submodules FIRST)
#############################
analyze -format sverilog ./${design_name}.sv

#############################
#  This assumes your top level module name is the file name without the extension
#############################
elaborate ${design_name}

#############################
#  Change this to match your clocks and timing constriaints
#############################
set_max_delay 25 -to [all_outputs]
create_clock "clk" -period 100
#create_clock "clk_in2" -period 100
#create_clock "clk_in3" -period 100

#############################
# if you have an internally generated clock instantiate a buffer (BUFX2)
# to provide a pin to identify the source of your new clock
#############################
#create_generated_clock -divide_by 1024 -source clk_in1 [get_pins {buffer/Y}]

report_clocks

check_design > check_design.output

ungroup -flatten -all

set_flatten true -effort high
uniquify

compile

#############################
# Check these files once completed 
#############################
report_area  > area.rpt
report_hierarchy > hierarchy.rpt
report_constraints > constraints.rpt
report_timing > timing.rpt

set_propagated_clock [all_clocks]

#############################
# Your timing file for IC Compiler 
#############################
write_sdc  ${design_name}.sdc

#############################
# Your output netlist 
#############################
write -f verilog ${design_name} -output ${design_name}.post_synth.v -hierarchy

# exit
                                                                                                                                                                                                                                                       adder_8.mag                                                                                         0000644 �    Asz0000145 00000004740 13045421026 010772  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1484427118
<< metal2 >>
rect 16 825 20 829
rect 8 809 12 813
rect 0 802 4 806
rect 16 715 20 820
rect 104 781 108 785
rect 8 699 12 703
rect 0 692 4 696
rect 16 605 20 710
rect 104 671 108 675
rect 8 589 12 593
rect 0 582 4 586
rect 16 495 20 600
rect 104 561 108 565
rect 8 479 12 483
rect 0 472 4 476
rect 16 385 20 490
rect 104 451 108 455
rect 8 369 12 373
rect 0 362 4 366
rect 16 275 20 380
rect 104 341 108 345
rect 8 259 12 263
rect 0 252 4 256
rect 16 165 20 270
rect 104 231 108 235
rect 8 149 12 153
rect 0 142 4 146
rect 16 55 20 162
rect 104 121 108 125
rect 16 47 20 51
rect 8 39 12 43
rect 0 32 4 36
rect 104 11 108 15
use fulladder  fulladder_0
timestamp 1484419411
transform 1 0 2 0 1 770
box -8 -4 128 96
use fulladder  fulladder_1
timestamp 1484419411
transform 1 0 2 0 1 660
box -8 -4 128 96
use fulladder  fulladder_2
timestamp 1484419411
transform 1 0 2 0 1 550
box -8 -4 128 96
use fulladder  fulladder_3
timestamp 1484419411
transform 1 0 2 0 1 440
box -8 -4 128 96
use fulladder  fulladder_4
timestamp 1484419411
transform 1 0 2 0 1 330
box -8 -4 128 96
use fulladder  fulladder_5
timestamp 1484419411
transform 1 0 2 0 1 220
box -8 -4 128 96
use fulladder  fulladder_6
timestamp 1484419411
transform 1 0 2 0 1 110
box -8 -4 128 96
use fulladder  fulladder_7
timestamp 1484419411
transform 1 0 2 0 1 0
box -8 -4 128 96
<< labels >>
rlabel metal2 1 34 1 34 1 a_0_
rlabel metal2 9 41 9 41 1 b_0_
rlabel metal2 1 144 1 144 1 a_1_
rlabel metal2 9 151 9 151 1 b_1_
rlabel metal2 0 252 4 256 1 a_2_
rlabel metal2 8 259 12 263 1 b_2_
rlabel metal2 0 362 4 366 1 a_3_
rlabel metal2 8 369 12 373 1 b_3_
rlabel metal2 0 472 4 476 1 a_4_
rlabel metal2 8 479 12 483 1 b_4_
rlabel metal2 0 582 4 586 1 a_5_
rlabel metal2 8 589 12 593 1 b_5_
rlabel metal2 0 692 4 696 1 a_6_
rlabel metal2 8 699 12 703 1 b_6_
rlabel metal2 0 802 4 806 1 a_7_
rlabel metal2 8 809 12 813 1 b_7_
rlabel metal2 16 47 20 51 1 cin
rlabel metal2 104 11 108 15 1 s_0_
rlabel metal2 104 121 108 125 1 s_1_
rlabel metal2 104 231 108 235 1 s_2_
rlabel metal2 104 341 108 345 1 s_3_
rlabel metal2 104 451 108 455 1 s_4_
rlabel metal2 104 561 108 565 1 s_5_
rlabel metal2 104 671 108 675 1 s_6_
rlabel metal2 104 781 108 785 1 s_7_
rlabel metal2 16 825 20 829 1 cout
rlabel metal2 16 715 20 719 1 c_7_
rlabel metal2 16 605 20 609 1 c_6_
rlabel metal2 16 495 20 499 1 c_5_
rlabel metal2 16 165 20 169 1 c_2_
rlabel metal2 16 55 20 59 1 c_1_
rlabel metal2 16 275 20 279 1 c_3_
rlabel metal2 16 385 20 389 1 c_4_
<< end >>
                                alt_alu.mag                                                                                         0000644 �    Asz0000145 00000001005 13050652047 011101  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1487098919
<< error_s >>
rect 29 157 36 159
use yzdetect_8  yzdetect_8_0
timestamp 1484534894
transform 1 0 8 0 1 4
box -8 -4 28 756
use inv_1x_8  inv_1x_8_0
timestamp 1484534894
transform 1 0 32 0 1 4
box -6 -4 18 866
use inv_1x_8  inv_1x_8_1
timestamp 1484534894
transform 1 0 48 0 1 4
box -6 -4 18 866
use adder_8  adder_8_0
timestamp 1484427118
transform 1 0 168 0 1 4
box -6 -4 130 866
use mux3_1x_8  mux3_1x_8_0
timestamp 1484532969
transform 1 0 296 0 1 4
box -6 -4 82 976
<< end >>
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           alt_alu_new.mag                                                                                     0000644 �    Asz0000145 00000040415 13055357611 011766  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1488314249
<< error_s >>
rect 84 100 92 101
<< nwell >>
rect 80 97 84 101
<< metal1 >>
rect 22 860 30 868
rect 22 770 30 778
rect 22 750 30 758
rect 22 660 30 668
rect 22 640 30 648
rect 22 550 30 558
rect 22 530 30 538
rect 22 440 30 448
rect 22 420 30 428
rect 22 330 30 338
rect 22 310 30 318
rect 22 220 30 228
rect 22 200 30 208
rect 22 110 30 118
rect 22 90 30 98
rect 22 0 30 8
<< m2contact >>
rect 352 763 356 767
<< metal2 >>
rect 184 926 188 927
rect 48 837 52 838
rect 32 824 33 827
rect 32 812 36 824
rect 40 806 44 816
rect 48 812 52 833
rect 144 837 148 838
rect 144 830 148 833
rect 184 833 188 922
rect 273 876 277 926
rect 296 922 300 938
rect 328 922 332 929
rect 56 819 60 820
rect 56 815 57 819
rect 56 812 60 815
rect 0 670 4 711
rect 16 690 20 776
rect 48 727 52 728
rect 32 714 33 717
rect 32 702 36 714
rect 40 696 44 706
rect 48 702 52 723
rect 56 709 60 710
rect 56 705 57 709
rect 56 702 60 705
rect 48 617 52 618
rect 32 604 33 607
rect 32 592 36 604
rect 40 586 44 596
rect 48 592 52 613
rect 56 599 60 600
rect 56 595 57 599
rect 56 592 60 595
rect 0 450 4 491
rect 23 474 27 556
rect 48 507 52 508
rect 32 494 33 497
rect 32 482 36 494
rect 40 476 44 486
rect 48 482 52 503
rect 56 489 60 490
rect 56 485 57 489
rect 56 482 60 485
rect 48 397 52 398
rect 32 384 33 387
rect 32 372 36 384
rect 8 367 12 371
rect 40 366 44 376
rect 48 372 52 393
rect 56 379 60 380
rect 56 375 57 379
rect 56 372 60 375
rect 0 230 4 271
rect 16 250 20 336
rect 48 287 52 288
rect 32 274 33 277
rect 32 262 36 274
rect 40 256 44 266
rect 48 262 52 283
rect 56 269 60 270
rect 56 265 57 269
rect 56 262 60 265
rect 48 177 52 178
rect 32 168 36 169
rect 32 152 36 164
rect 40 146 44 156
rect 48 152 52 173
rect 56 159 60 160
rect 56 155 57 159
rect 56 152 60 155
rect 0 10 4 51
rect 16 30 20 116
rect 80 101 84 812
rect 48 67 52 68
rect 32 54 33 57
rect 32 42 36 54
rect 40 36 44 46
rect 48 42 52 63
rect 56 49 60 50
rect 56 45 57 49
rect 56 42 60 45
rect 80 38 84 97
rect 88 321 92 812
rect 112 806 116 812
rect 112 696 116 702
rect 112 586 116 592
rect 120 541 124 827
rect 160 811 164 813
rect 112 476 116 482
rect 112 366 116 372
rect 88 38 92 317
rect 112 256 116 262
rect 112 146 116 152
rect 96 53 100 54
rect 120 53 124 537
rect 136 761 140 811
rect 168 806 172 824
rect 312 817 316 826
rect 304 789 308 817
rect 112 36 116 42
rect 136 37 140 757
rect 144 727 148 728
rect 144 720 148 723
rect 160 701 164 703
rect 168 696 172 714
rect 312 707 316 716
rect 304 679 308 707
rect 144 617 148 618
rect 144 610 148 613
rect 160 591 164 593
rect 168 586 172 604
rect 312 597 316 606
rect 304 569 308 597
rect 144 507 148 508
rect 144 500 148 503
rect 160 481 164 483
rect 168 476 172 494
rect 312 487 316 496
rect 304 459 308 487
rect 144 397 148 398
rect 144 390 148 393
rect 160 371 164 373
rect 168 366 172 384
rect 312 377 316 386
rect 304 349 308 377
rect 144 287 148 288
rect 144 280 148 283
rect 160 261 164 263
rect 168 256 172 274
rect 312 267 316 276
rect 304 239 308 267
rect 144 177 148 178
rect 144 170 148 173
rect 160 151 164 153
rect 168 146 172 164
rect 312 157 316 166
rect 304 129 308 157
rect 144 67 148 68
rect 144 60 148 63
rect 279 58 283 106
rect 160 41 164 43
rect 168 36 172 54
rect 328 56 332 872
rect 352 767 356 826
rect 368 780 372 816
rect 352 104 356 763
rect 379 761 383 763
rect 368 670 372 706
rect 379 702 383 757
rect 368 560 372 596
rect 379 492 383 537
rect 368 450 372 486
rect 368 340 372 376
rect 379 272 383 317
rect 368 230 372 266
rect 368 120 372 156
rect 389 110 393 917
rect 379 62 383 97
rect 184 51 188 52
rect 312 47 316 56
rect 304 19 308 47
rect 368 10 372 46
<< m3contact >>
rect 296 938 300 942
rect 691 938 695 942
rect 184 922 188 926
rect 265 922 269 926
rect 48 833 52 837
rect 33 824 37 828
rect 144 833 148 837
rect 328 929 332 933
rect 395 929 399 933
rect 389 917 393 921
rect 273 872 277 876
rect 328 872 332 876
rect 184 829 188 833
rect 95 824 100 828
rect 57 815 61 819
rect 64 815 68 819
rect 40 802 44 806
rect 16 776 20 780
rect 48 723 52 727
rect 33 714 37 718
rect 57 705 61 709
rect 64 705 68 709
rect 40 692 44 696
rect 0 666 4 670
rect 48 613 52 617
rect 33 604 37 608
rect 57 595 61 599
rect 64 595 68 599
rect 40 582 44 586
rect 23 556 27 560
rect 48 503 52 507
rect 33 494 37 498
rect 16 470 20 474
rect 23 470 27 474
rect 57 485 61 489
rect 64 485 68 489
rect 40 472 44 476
rect 0 446 4 450
rect 48 393 52 397
rect 33 384 37 388
rect 57 375 61 379
rect 64 375 68 379
rect 40 362 44 366
rect 16 336 20 340
rect 48 283 52 287
rect 33 274 37 278
rect 57 265 61 269
rect 64 265 68 269
rect 40 252 44 256
rect 0 226 4 230
rect 48 173 52 177
rect 32 164 36 168
rect 57 155 61 159
rect 64 155 68 159
rect 40 142 44 146
rect 16 116 20 120
rect 80 97 84 101
rect 48 63 52 67
rect 33 54 37 58
rect 57 45 61 49
rect 64 45 68 49
rect 112 802 116 806
rect 95 714 100 718
rect 112 692 116 696
rect 95 604 100 608
rect 112 582 116 586
rect 168 824 172 828
rect 160 813 164 817
rect 120 537 124 541
rect 95 494 100 498
rect 112 472 116 476
rect 95 384 100 388
rect 112 362 116 366
rect 88 317 92 321
rect 95 274 100 278
rect 112 252 116 256
rect 95 164 100 168
rect 112 142 116 146
rect 95 54 100 58
rect 176 813 180 817
rect 312 813 316 817
rect 272 785 276 789
rect 304 785 308 789
rect 136 757 140 761
rect 40 32 44 36
rect 144 723 148 727
rect 168 714 172 718
rect 160 703 164 707
rect 176 703 180 707
rect 312 703 316 707
rect 272 675 276 679
rect 304 675 308 679
rect 144 613 148 617
rect 168 604 172 608
rect 160 593 164 597
rect 176 593 180 597
rect 312 593 316 597
rect 272 565 276 569
rect 304 565 308 569
rect 144 503 148 507
rect 168 494 172 498
rect 160 483 164 487
rect 176 483 180 487
rect 312 483 316 487
rect 272 455 276 459
rect 304 455 308 459
rect 144 393 148 397
rect 168 384 172 388
rect 160 373 164 377
rect 176 373 180 377
rect 312 373 316 377
rect 272 345 276 349
rect 304 345 308 349
rect 144 283 148 287
rect 168 274 172 278
rect 160 263 164 267
rect 176 263 180 267
rect 312 263 316 267
rect 272 235 276 239
rect 304 235 308 239
rect 144 173 148 177
rect 168 164 172 168
rect 160 153 164 157
rect 176 153 180 157
rect 312 153 316 157
rect 272 125 276 129
rect 304 125 308 129
rect 279 106 283 110
rect 144 63 148 67
rect 168 54 172 58
rect 160 43 164 47
rect 184 52 188 56
rect 279 54 283 58
rect 368 776 372 780
rect 379 757 383 761
rect 379 698 383 702
rect 368 666 372 670
rect 368 556 372 560
rect 379 537 383 541
rect 379 488 383 492
rect 368 446 372 450
rect 368 336 372 340
rect 379 317 383 321
rect 379 268 383 272
rect 368 226 372 230
rect 368 116 372 120
rect 389 106 393 110
rect 379 97 383 101
rect 379 58 383 62
rect 328 52 332 56
rect 352 52 356 56
rect 176 43 180 47
rect 112 32 116 36
rect 312 43 316 47
rect 272 15 276 19
rect 304 15 308 19
rect 0 6 4 10
rect 368 6 372 10
<< metal3 >>
rect 295 942 697 943
rect 295 938 296 942
rect 300 938 691 942
rect 695 938 697 942
rect 295 937 697 938
rect 327 933 400 934
rect 327 929 328 933
rect 332 929 395 933
rect 399 929 400 933
rect 327 928 400 929
rect 183 926 270 927
rect 183 922 184 926
rect 188 922 265 926
rect 269 922 270 926
rect 183 921 270 922
rect 388 921 394 922
rect 388 917 389 921
rect 393 917 394 921
rect 388 916 394 917
rect 272 876 333 877
rect 272 872 273 876
rect 277 872 328 876
rect 332 872 333 876
rect 272 871 333 872
rect 47 837 149 838
rect 47 833 48 837
rect 52 833 144 837
rect 148 833 149 837
rect 47 832 149 833
rect 183 833 189 834
rect 183 829 184 833
rect 188 829 189 833
rect 32 828 173 829
rect 183 828 189 829
rect 32 824 33 828
rect 37 824 95 828
rect 100 824 168 828
rect 172 824 173 828
rect 32 823 173 824
rect 56 819 69 820
rect 56 815 57 819
rect 61 815 64 819
rect 68 815 69 819
rect 56 814 69 815
rect 159 817 317 818
rect 159 813 160 817
rect 164 813 176 817
rect 180 813 312 817
rect 316 813 317 817
rect 159 812 317 813
rect 39 806 117 807
rect 39 802 40 806
rect 44 802 112 806
rect 116 802 117 806
rect 39 801 117 802
rect 271 789 309 790
rect 271 785 272 789
rect 276 785 304 789
rect 308 785 309 789
rect 271 784 309 785
rect -2 780 373 781
rect -2 776 16 780
rect 20 776 368 780
rect 372 776 373 780
rect -2 775 373 776
rect 135 761 384 762
rect 135 757 136 761
rect 140 757 379 761
rect 383 757 384 761
rect 135 756 384 757
rect 47 727 149 728
rect 47 723 48 727
rect 52 723 144 727
rect 148 723 149 727
rect 47 722 149 723
rect 32 718 173 719
rect 32 714 33 718
rect 37 714 95 718
rect 100 714 168 718
rect 172 714 173 718
rect 32 713 173 714
rect 56 709 69 710
rect 56 705 57 709
rect 61 705 64 709
rect 68 705 69 709
rect 56 704 69 705
rect 159 707 317 708
rect 159 703 160 707
rect 164 703 176 707
rect 180 703 312 707
rect 316 703 317 707
rect 159 702 317 703
rect 378 702 384 703
rect 378 698 379 702
rect 383 698 384 702
rect 378 697 384 698
rect 39 696 117 697
rect 39 692 40 696
rect 44 692 112 696
rect 116 692 117 696
rect 39 691 117 692
rect 271 679 309 680
rect 271 675 272 679
rect 276 675 304 679
rect 308 675 309 679
rect 271 674 309 675
rect -2 670 373 671
rect -2 666 0 670
rect 4 666 368 670
rect 372 666 373 670
rect -2 665 373 666
rect 47 617 149 618
rect 47 613 48 617
rect 52 613 144 617
rect 148 613 149 617
rect 47 612 149 613
rect 32 608 173 609
rect 32 604 33 608
rect 37 604 95 608
rect 100 604 168 608
rect 172 604 173 608
rect 32 603 173 604
rect 56 599 69 600
rect 56 595 57 599
rect 61 595 64 599
rect 68 595 69 599
rect 56 594 69 595
rect 159 597 317 598
rect 159 593 160 597
rect 164 593 176 597
rect 180 593 312 597
rect 316 593 317 597
rect 159 592 317 593
rect 39 586 117 587
rect 39 582 40 586
rect 44 582 112 586
rect 116 582 117 586
rect 39 581 117 582
rect 271 569 309 570
rect 271 565 272 569
rect 276 565 304 569
rect 308 565 309 569
rect 271 564 309 565
rect -2 560 373 561
rect -2 556 23 560
rect 27 556 368 560
rect 372 556 373 560
rect -2 555 373 556
rect 119 541 384 542
rect 119 537 120 541
rect 124 537 379 541
rect 383 537 384 541
rect 119 536 384 537
rect 47 507 149 508
rect 47 503 48 507
rect 52 503 144 507
rect 148 503 149 507
rect 47 502 149 503
rect 32 498 173 499
rect 32 494 33 498
rect 37 494 95 498
rect 100 494 168 498
rect 172 494 173 498
rect 32 493 173 494
rect 378 492 384 493
rect 56 489 69 490
rect 56 485 57 489
rect 61 485 64 489
rect 68 485 69 489
rect 378 488 379 492
rect 383 488 384 492
rect 56 484 69 485
rect 159 487 317 488
rect 378 487 384 488
rect 159 483 160 487
rect 164 483 176 487
rect 180 483 312 487
rect 316 483 317 487
rect 159 482 317 483
rect 39 476 117 477
rect 15 474 28 475
rect 15 470 16 474
rect 20 470 23 474
rect 27 470 28 474
rect 39 472 40 476
rect 44 472 112 476
rect 116 472 117 476
rect 39 471 117 472
rect 15 469 28 470
rect 271 459 309 460
rect 271 455 272 459
rect 276 455 304 459
rect 308 455 309 459
rect 271 454 309 455
rect -2 450 373 451
rect -2 446 0 450
rect 4 446 368 450
rect 372 446 373 450
rect -2 445 373 446
rect 47 397 149 398
rect 47 393 48 397
rect 52 393 144 397
rect 148 393 149 397
rect 47 392 149 393
rect 32 388 173 389
rect 32 384 33 388
rect 37 384 95 388
rect 100 384 168 388
rect 172 384 173 388
rect 32 383 173 384
rect 56 379 69 380
rect 56 375 57 379
rect 61 375 64 379
rect 68 375 69 379
rect 56 374 69 375
rect 159 377 317 378
rect 159 373 160 377
rect 164 373 176 377
rect 180 373 312 377
rect 316 373 317 377
rect 159 372 317 373
rect 39 366 117 367
rect 39 362 40 366
rect 44 362 112 366
rect 116 362 117 366
rect 39 361 117 362
rect 271 349 309 350
rect 271 345 272 349
rect 276 345 304 349
rect 308 345 309 349
rect 271 344 309 345
rect -2 340 373 341
rect -2 336 16 340
rect 20 336 368 340
rect 372 336 373 340
rect -2 335 373 336
rect 87 321 384 322
rect 87 317 88 321
rect 92 317 379 321
rect 383 317 384 321
rect 87 316 384 317
rect 47 287 149 288
rect 47 283 48 287
rect 52 283 144 287
rect 148 283 149 287
rect 47 282 149 283
rect 32 278 173 279
rect 32 274 33 278
rect 37 274 95 278
rect 100 274 168 278
rect 172 274 173 278
rect 32 273 173 274
rect 378 272 384 273
rect 56 269 69 270
rect 56 265 57 269
rect 61 265 64 269
rect 68 265 69 269
rect 378 268 379 272
rect 383 268 384 272
rect 56 264 69 265
rect 159 267 317 268
rect 378 267 384 268
rect 159 263 160 267
rect 164 263 176 267
rect 180 263 312 267
rect 316 263 317 267
rect 159 262 317 263
rect 39 256 117 257
rect 39 252 40 256
rect 44 252 112 256
rect 116 252 117 256
rect 39 251 117 252
rect 271 239 309 240
rect 271 235 272 239
rect 276 235 304 239
rect 308 235 309 239
rect 271 234 309 235
rect -2 230 373 231
rect -2 226 0 230
rect 4 226 368 230
rect 372 226 373 230
rect -2 225 373 226
rect 47 177 149 178
rect 47 173 48 177
rect 52 173 144 177
rect 148 173 149 177
rect 47 172 149 173
rect 31 168 173 169
rect 31 164 32 168
rect 36 164 95 168
rect 100 164 168 168
rect 172 164 173 168
rect 31 163 173 164
rect 56 159 69 160
rect 56 155 57 159
rect 61 155 64 159
rect 68 155 69 159
rect 56 154 69 155
rect 159 157 317 158
rect 159 153 160 157
rect 164 153 176 157
rect 180 153 312 157
rect 316 153 317 157
rect 159 152 317 153
rect 39 146 117 147
rect 39 142 40 146
rect 44 142 112 146
rect 116 142 117 146
rect 39 141 117 142
rect 271 129 309 130
rect 271 125 272 129
rect 276 125 304 129
rect 308 125 309 129
rect 271 124 309 125
rect -2 120 373 121
rect -2 116 16 120
rect 20 116 368 120
rect 372 116 373 120
rect -2 115 373 116
rect 278 110 395 111
rect 278 106 279 110
rect 283 106 389 110
rect 393 106 395 110
rect 278 105 395 106
rect 79 101 384 102
rect 79 97 80 101
rect 84 97 379 101
rect 383 97 384 101
rect 79 96 384 97
rect 47 67 149 68
rect 47 63 48 67
rect 52 63 144 67
rect 148 63 149 67
rect 47 62 149 63
rect 378 62 384 63
rect 32 58 173 59
rect 32 54 33 58
rect 37 54 95 58
rect 100 54 168 58
rect 172 54 173 58
rect 32 53 173 54
rect 183 58 284 59
rect 183 56 279 58
rect 183 52 184 56
rect 188 54 279 56
rect 283 54 284 58
rect 378 58 379 62
rect 383 58 384 62
rect 378 57 384 58
rect 188 53 284 54
rect 327 56 357 57
rect 188 52 189 53
rect 183 51 189 52
rect 327 52 328 56
rect 332 52 352 56
rect 356 52 357 56
rect 327 51 357 52
rect 56 49 69 50
rect 56 45 57 49
rect 61 45 64 49
rect 68 45 69 49
rect 56 44 69 45
rect 159 47 317 48
rect 159 43 160 47
rect 164 43 176 47
rect 180 43 312 47
rect 316 43 317 47
rect 159 42 317 43
rect 39 36 117 37
rect 39 32 40 36
rect 44 32 112 36
rect 116 32 117 36
rect 39 31 117 32
rect 271 19 309 20
rect 271 15 272 19
rect 276 15 304 19
rect 308 15 309 19
rect 271 14 309 15
rect -2 10 373 11
rect -2 6 0 10
rect 4 6 368 10
rect 372 6 373 10
rect -2 5 373 6
use inv_1x  inv_1x_0
timestamp 1484418501
transform 1 0 265 0 1 884
box -6 -4 18 96
use yzdetect_8  yzdetect_8_0
timestamp 1484534894
transform 1 0 0 0 1 4
box -8 -4 28 756
use inv_1x_8  inv_1x_8_0
timestamp 1484534894
transform 1 0 32 0 1 4
box -6 -4 18 866
use inv_1x_8  inv_1x_8_1
timestamp 1484534894
transform 1 0 48 0 1 4
box -6 -4 18 866
use mux4_8_10space  mux4_8_10space_0
timestamp 1487099744
transform 1 0 58 0 1 0
box 0 0 112 870
use adder_8  adder_8_0
timestamp 1484427118
transform 1 0 168 0 1 4
box -6 -4 130 866
use mux3_1x_8  mux3_1x_8_0
timestamp 1484532969
transform 1 0 296 0 1 4
box -6 -4 82 976
use alu_ctl  alu_ctl_0
timestamp 1488311641
transform 1 0 378 0 1 0
box 0 0 400 980
<< labels >>
rlabel metal2 33 46 33 46 1 a0
rlabel metal2 49 46 49 46 1 b0
rlabel metal2 33 156 33 156 1 a1
rlabel metal2 49 156 49 156 1 b1
rlabel metal2 33 266 33 266 1 a2
rlabel metal2 49 266 49 266 1 b2
rlabel metal2 33 376 33 376 1 a3
rlabel metal2 49 376 49 376 1 b3
rlabel metal2 33 486 33 486 1 a4
rlabel metal2 49 486 49 486 1 b4
rlabel metal2 33 596 33 596 1 a5
rlabel metal3 -1 9 -1 9 1 result0
rlabel metal3 -1 119 -1 119 1 result1
rlabel metal3 -1 230 -1 230 1 result2
rlabel metal3 -1 340 -1 340 1 result3
rlabel metal3 -1 450 -1 450 1 result4
rlabel metal3 -1 560 -1 560 1 result5
rlabel metal3 -1 670 -1 670 1 result6
rlabel metal3 1 778 1 778 1 result7
rlabel m2contact 352 763 356 767 1 less
rlabel metal2 296 922 300 926 1 op0
rlabel metal2 328 922 332 926 1 op1
rlabel metal2 49 596 49 596 1 b5
rlabel metal2 33 706 33 706 1 a6
rlabel metal2 49 706 49 706 1 b6
rlabel metal2 33 816 33 816 1 a7
rlabel metal2 49 816 49 816 1 b7
rlabel metal2 9 370 9 370 1 zero
rlabel m3contact 161 44 161 44 1 muxy7
rlabel metal2 81 767 81 767 1 op6
rlabel metal2 89 767 89 767 1 op5
rlabel metal2 120 763 124 767 1 op4
rlabel metal2 136 763 140 767 1 op3
rlabel m3contact 98 56 98 56 1 mux4s1_0
rlabel metal2 146 61 146 61 1 mux4s0_0
rlabel m3contact 186 830 186 830 1 cout_adder_7
rlabel metal2 122 544 122 544 1 op4
rlabel metal2 90 325 90 325 1 op5
rlabel metal2 82 104 82 104 1 op6
rlabel metal2 186 52 186 52 1 op2
rlabel metal2 281 106 281 106 1 op2
<< end >>
                                                                                                                                                                                                                                                   alt_alu_with_ctl.mag                                                                                0000644 �    Asz0000145 00000043120 13055370460 013003  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1488318768
<< metal1 >>
rect 22 860 30 868
rect 22 770 30 778
rect 22 750 30 758
rect 22 660 30 668
rect 22 640 30 648
rect 22 550 30 558
rect 22 530 30 538
rect 22 440 30 448
rect 22 420 30 428
rect 22 330 30 338
rect 22 310 30 318
rect 22 220 30 228
rect 22 200 30 208
rect 22 110 30 118
rect 22 90 30 98
rect 22 0 30 8
<< m2contact >>
rect 352 763 356 767
rect 555 69 559 73
rect 552 43 556 47
<< metal2 >>
rect 184 926 188 927
rect 48 837 52 838
rect 32 824 33 827
rect 32 812 36 824
rect 40 806 44 816
rect 48 812 52 833
rect 144 837 148 838
rect 144 830 148 833
rect 184 833 188 922
rect 273 876 277 926
rect 296 922 300 938
rect 328 922 332 929
rect 770 918 771 922
rect 775 918 778 922
rect 770 917 778 918
rect 56 819 60 820
rect 56 815 57 819
rect 56 812 60 815
rect 0 670 4 711
rect 16 690 20 776
rect 48 727 52 728
rect 32 714 33 717
rect 32 702 36 714
rect 40 696 44 706
rect 48 702 52 723
rect 56 709 60 710
rect 56 705 57 709
rect 56 702 60 705
rect 48 617 52 618
rect 32 604 33 607
rect 32 592 36 604
rect 40 586 44 596
rect 48 592 52 613
rect 56 599 60 600
rect 56 595 57 599
rect 56 592 60 595
rect 0 450 4 491
rect 23 474 27 556
rect 48 507 52 508
rect 32 494 33 497
rect 32 482 36 494
rect 40 476 44 486
rect 48 482 52 503
rect 56 489 60 490
rect 56 485 57 489
rect 56 482 60 485
rect 48 397 52 398
rect 32 384 33 387
rect 32 372 36 384
rect 8 367 12 371
rect 40 366 44 376
rect 48 372 52 393
rect 56 379 60 380
rect 56 375 57 379
rect 56 372 60 375
rect 0 230 4 271
rect 16 250 20 336
rect 48 287 52 288
rect 32 274 33 277
rect 32 262 36 274
rect 40 256 44 266
rect 48 262 52 283
rect 56 269 60 270
rect 56 265 57 269
rect 56 262 60 265
rect 48 177 52 178
rect 32 168 36 169
rect 32 152 36 164
rect 40 146 44 156
rect 48 152 52 173
rect 56 159 60 160
rect 56 155 57 159
rect 56 152 60 155
rect 0 10 4 51
rect 16 30 20 116
rect 80 101 84 812
rect 48 67 52 68
rect 32 54 33 57
rect 32 42 36 54
rect 40 36 44 46
rect 48 42 52 63
rect 56 49 60 50
rect 56 45 57 49
rect 56 42 60 45
rect 80 38 84 97
rect 88 321 92 812
rect 112 806 116 812
rect 112 696 116 702
rect 112 586 116 592
rect 120 541 124 827
rect 160 811 164 813
rect 112 476 116 482
rect 112 366 116 372
rect 88 38 92 317
rect 112 256 116 262
rect 112 146 116 152
rect 96 53 100 54
rect 120 53 124 537
rect 136 761 140 811
rect 168 806 172 824
rect 312 817 316 826
rect 304 789 308 817
rect 112 36 116 42
rect 136 37 140 757
rect 144 727 148 728
rect 144 720 148 723
rect 160 701 164 703
rect 168 696 172 714
rect 312 707 316 716
rect 304 679 308 707
rect 144 617 148 618
rect 144 610 148 613
rect 160 591 164 593
rect 168 586 172 604
rect 312 597 316 606
rect 304 569 308 597
rect 144 507 148 508
rect 144 500 148 503
rect 160 481 164 483
rect 168 476 172 494
rect 312 487 316 496
rect 304 459 308 487
rect 144 397 148 398
rect 144 390 148 393
rect 160 371 164 373
rect 168 366 172 384
rect 312 377 316 386
rect 304 349 308 377
rect 144 287 148 288
rect 144 280 148 283
rect 160 261 164 263
rect 168 256 172 274
rect 312 267 316 276
rect 304 239 308 267
rect 144 177 148 178
rect 144 170 148 173
rect 160 151 164 153
rect 168 146 172 164
rect 312 157 316 166
rect 304 129 308 157
rect 144 67 148 68
rect 144 60 148 63
rect 279 58 283 106
rect 160 41 164 43
rect 168 36 172 54
rect 328 56 332 872
rect 352 767 356 826
rect 368 780 372 816
rect 352 104 356 763
rect 379 761 383 763
rect 368 670 372 706
rect 379 702 383 757
rect 368 560 372 596
rect 379 492 383 537
rect 368 450 372 486
rect 368 340 372 376
rect 379 272 383 317
rect 368 230 372 266
rect 368 120 372 156
rect 389 110 393 917
rect 768 698 769 702
rect 773 698 776 702
rect 768 697 776 698
rect 769 488 770 492
rect 774 488 777 492
rect 769 487 777 488
rect 766 268 770 272
rect 774 268 778 272
rect 766 267 778 268
rect 379 62 383 97
rect 768 61 776 62
rect 768 57 769 61
rect 773 57 776 61
rect 184 51 188 52
rect 312 47 316 56
rect 304 19 308 47
rect 368 10 372 46
rect 404 0 412 3
rect 716 0 723 3
<< m3contact >>
rect 296 938 300 942
rect 691 938 695 942
rect 184 922 188 926
rect 265 922 269 926
rect 48 833 52 837
rect 33 824 37 828
rect 144 833 148 837
rect 328 929 332 933
rect 395 929 399 933
rect 389 917 393 921
rect 771 918 775 922
rect 273 872 277 876
rect 328 872 332 876
rect 184 829 188 833
rect 95 824 100 828
rect 57 815 61 819
rect 64 815 68 819
rect 40 802 44 806
rect 16 776 20 780
rect 48 723 52 727
rect 33 714 37 718
rect 57 705 61 709
rect 64 705 68 709
rect 40 692 44 696
rect 0 666 4 670
rect 48 613 52 617
rect 33 604 37 608
rect 57 595 61 599
rect 64 595 68 599
rect 40 582 44 586
rect 23 556 27 560
rect 48 503 52 507
rect 33 494 37 498
rect 16 470 20 474
rect 23 470 27 474
rect 57 485 61 489
rect 64 485 68 489
rect 40 472 44 476
rect 0 446 4 450
rect 48 393 52 397
rect 33 384 37 388
rect 57 375 61 379
rect 64 375 68 379
rect 40 362 44 366
rect 16 336 20 340
rect 48 283 52 287
rect 33 274 37 278
rect 57 265 61 269
rect 64 265 68 269
rect 40 252 44 256
rect 0 226 4 230
rect 48 173 52 177
rect 32 164 36 168
rect 57 155 61 159
rect 64 155 68 159
rect 40 142 44 146
rect 16 116 20 120
rect 80 97 84 101
rect 48 63 52 67
rect 33 54 37 58
rect 57 45 61 49
rect 64 45 68 49
rect 112 802 116 806
rect 95 714 100 718
rect 112 692 116 696
rect 95 604 100 608
rect 112 582 116 586
rect 168 824 172 828
rect 160 813 164 817
rect 120 537 124 541
rect 95 494 100 498
rect 112 472 116 476
rect 95 384 100 388
rect 112 362 116 366
rect 88 317 92 321
rect 95 274 100 278
rect 112 252 116 256
rect 95 164 100 168
rect 112 142 116 146
rect 95 54 100 58
rect 176 813 180 817
rect 312 813 316 817
rect 272 785 276 789
rect 304 785 308 789
rect 136 757 140 761
rect 40 32 44 36
rect 144 723 148 727
rect 168 714 172 718
rect 160 703 164 707
rect 176 703 180 707
rect 312 703 316 707
rect 272 675 276 679
rect 304 675 308 679
rect 144 613 148 617
rect 168 604 172 608
rect 160 593 164 597
rect 176 593 180 597
rect 312 593 316 597
rect 272 565 276 569
rect 304 565 308 569
rect 144 503 148 507
rect 168 494 172 498
rect 160 483 164 487
rect 176 483 180 487
rect 312 483 316 487
rect 272 455 276 459
rect 304 455 308 459
rect 144 393 148 397
rect 168 384 172 388
rect 160 373 164 377
rect 176 373 180 377
rect 312 373 316 377
rect 272 345 276 349
rect 304 345 308 349
rect 144 283 148 287
rect 168 274 172 278
rect 160 263 164 267
rect 176 263 180 267
rect 312 263 316 267
rect 272 235 276 239
rect 304 235 308 239
rect 144 173 148 177
rect 168 164 172 168
rect 160 153 164 157
rect 176 153 180 157
rect 312 153 316 157
rect 272 125 276 129
rect 304 125 308 129
rect 279 106 283 110
rect 144 63 148 67
rect 168 54 172 58
rect 160 43 164 47
rect 184 52 188 56
rect 279 54 283 58
rect 368 776 372 780
rect 379 757 383 761
rect 379 698 383 702
rect 368 666 372 670
rect 368 556 372 560
rect 379 537 383 541
rect 379 488 383 492
rect 379 468 383 472
rect 368 446 372 450
rect 368 336 372 340
rect 379 317 383 321
rect 379 268 383 272
rect 368 226 372 230
rect 368 116 372 120
rect 769 698 773 702
rect 770 488 774 492
rect 770 268 774 272
rect 389 106 393 110
rect 379 97 383 101
rect 379 58 383 62
rect 769 57 773 61
rect 328 52 332 56
rect 352 52 356 56
rect 176 43 180 47
rect 112 32 116 36
rect 312 43 316 47
rect 272 15 276 19
rect 304 15 308 19
rect 0 6 4 10
rect 368 6 372 10
<< metal3 >>
rect 295 942 697 943
rect 295 938 296 942
rect 300 938 691 942
rect 695 938 697 942
rect 295 937 697 938
rect 327 933 400 934
rect 327 929 328 933
rect 332 929 395 933
rect 399 929 400 933
rect 327 928 400 929
rect 183 926 270 927
rect 183 922 184 926
rect 188 922 265 926
rect 269 922 270 926
rect 770 922 776 923
rect 183 921 270 922
rect 388 921 394 922
rect 388 917 389 921
rect 393 917 394 921
rect 770 918 771 922
rect 775 918 778 922
rect 770 917 778 918
rect 388 916 394 917
rect 272 876 333 877
rect 272 872 273 876
rect 277 872 328 876
rect 332 872 333 876
rect 272 871 333 872
rect 47 837 149 838
rect 47 833 48 837
rect 52 833 144 837
rect 148 833 149 837
rect 47 832 149 833
rect 183 833 189 834
rect 183 829 184 833
rect 188 829 189 833
rect 32 828 173 829
rect 183 828 189 829
rect 32 824 33 828
rect 37 824 95 828
rect 100 824 168 828
rect 172 824 173 828
rect 32 823 173 824
rect 56 819 69 820
rect 56 815 57 819
rect 61 815 64 819
rect 68 815 69 819
rect 56 814 69 815
rect 159 817 317 818
rect 159 813 160 817
rect 164 813 176 817
rect 180 813 312 817
rect 316 813 317 817
rect 159 812 317 813
rect 39 806 117 807
rect 39 802 40 806
rect 44 802 112 806
rect 116 802 117 806
rect 39 801 117 802
rect 271 789 309 790
rect 271 785 272 789
rect 276 785 304 789
rect 308 785 309 789
rect 271 784 309 785
rect -2 780 373 781
rect -2 776 16 780
rect 20 776 368 780
rect 372 776 373 780
rect -2 775 373 776
rect 135 761 384 762
rect 135 757 136 761
rect 140 757 379 761
rect 383 757 384 761
rect 135 756 384 757
rect 47 727 149 728
rect 47 723 48 727
rect 52 723 144 727
rect 148 723 149 727
rect 47 722 149 723
rect 32 718 173 719
rect 32 714 33 718
rect 37 714 95 718
rect 100 714 168 718
rect 172 714 173 718
rect 32 713 173 714
rect 56 709 69 710
rect 56 705 57 709
rect 61 705 64 709
rect 68 705 69 709
rect 56 704 69 705
rect 159 707 317 708
rect 159 703 160 707
rect 164 703 176 707
rect 180 703 312 707
rect 316 703 317 707
rect 159 702 317 703
rect 378 702 384 703
rect 378 698 379 702
rect 383 698 384 702
rect 378 697 384 698
rect 768 702 774 703
rect 768 698 769 702
rect 773 698 776 702
rect 768 697 776 698
rect 39 696 117 697
rect 39 692 40 696
rect 44 692 112 696
rect 116 692 117 696
rect 39 691 117 692
rect 271 679 309 680
rect 271 675 272 679
rect 276 675 304 679
rect 308 675 309 679
rect 271 674 309 675
rect -2 670 373 671
rect -2 666 0 670
rect 4 666 368 670
rect 372 666 373 670
rect -2 665 373 666
rect 47 617 149 618
rect 47 613 48 617
rect 52 613 144 617
rect 148 613 149 617
rect 47 612 149 613
rect 32 608 173 609
rect 32 604 33 608
rect 37 604 95 608
rect 100 604 168 608
rect 172 604 173 608
rect 32 603 173 604
rect 56 599 69 600
rect 56 595 57 599
rect 61 595 64 599
rect 68 595 69 599
rect 56 594 69 595
rect 159 597 317 598
rect 159 593 160 597
rect 164 593 176 597
rect 180 593 312 597
rect 316 593 317 597
rect 159 592 317 593
rect 39 586 117 587
rect 39 582 40 586
rect 44 582 112 586
rect 116 582 117 586
rect 39 581 117 582
rect 271 569 309 570
rect 271 565 272 569
rect 276 565 304 569
rect 308 565 309 569
rect 271 564 309 565
rect -2 560 373 561
rect -2 556 23 560
rect 27 556 368 560
rect 372 556 373 560
rect -2 555 373 556
rect 119 541 384 542
rect 119 537 120 541
rect 124 537 379 541
rect 383 537 384 541
rect 119 536 384 537
rect 47 507 149 508
rect 47 503 48 507
rect 52 503 144 507
rect 148 503 149 507
rect 47 502 149 503
rect 32 498 173 499
rect 32 494 33 498
rect 37 494 95 498
rect 100 494 168 498
rect 172 494 173 498
rect 32 493 173 494
rect 378 492 384 493
rect 56 489 69 490
rect 56 485 57 489
rect 61 485 64 489
rect 68 485 69 489
rect 378 488 379 492
rect 383 488 384 492
rect 56 484 69 485
rect 159 487 317 488
rect 378 487 384 488
rect 769 492 775 493
rect 769 488 770 492
rect 774 488 777 492
rect 769 487 777 488
rect 159 483 160 487
rect 164 483 176 487
rect 180 483 312 487
rect 316 483 317 487
rect 159 482 317 483
rect 39 476 117 477
rect 15 474 28 475
rect 15 470 16 474
rect 20 470 23 474
rect 27 470 28 474
rect 39 472 40 476
rect 44 472 112 476
rect 116 472 117 476
rect 39 471 117 472
rect 378 472 384 473
rect 15 469 28 470
rect 378 468 379 472
rect 383 468 384 472
rect 378 467 384 468
rect 271 459 309 460
rect 271 455 272 459
rect 276 455 304 459
rect 308 455 309 459
rect 271 454 309 455
rect -2 450 373 451
rect -2 446 0 450
rect 4 446 368 450
rect 372 446 373 450
rect -2 445 373 446
rect 47 397 149 398
rect 47 393 48 397
rect 52 393 144 397
rect 148 393 149 397
rect 47 392 149 393
rect 32 388 173 389
rect 32 384 33 388
rect 37 384 95 388
rect 100 384 168 388
rect 172 384 173 388
rect 32 383 173 384
rect 56 379 69 380
rect 56 375 57 379
rect 61 375 64 379
rect 68 375 69 379
rect 56 374 69 375
rect 159 377 317 378
rect 159 373 160 377
rect 164 373 176 377
rect 180 373 312 377
rect 316 373 317 377
rect 159 372 317 373
rect 39 366 117 367
rect 39 362 40 366
rect 44 362 112 366
rect 116 362 117 366
rect 39 361 117 362
rect 271 349 309 350
rect 271 345 272 349
rect 276 345 304 349
rect 308 345 309 349
rect 271 344 309 345
rect -2 340 373 341
rect -2 336 16 340
rect 20 336 368 340
rect 372 336 373 340
rect -2 335 373 336
rect 87 321 384 322
rect 87 317 88 321
rect 92 317 379 321
rect 383 317 384 321
rect 87 316 384 317
rect 47 287 149 288
rect 47 283 48 287
rect 52 283 144 287
rect 148 283 149 287
rect 47 282 149 283
rect 32 278 173 279
rect 32 274 33 278
rect 37 274 95 278
rect 100 274 168 278
rect 172 274 173 278
rect 32 273 173 274
rect 378 272 384 273
rect 769 272 775 273
rect 56 269 69 270
rect 56 265 57 269
rect 61 265 64 269
rect 68 265 69 269
rect 378 268 379 272
rect 383 268 384 272
rect 56 264 69 265
rect 159 267 317 268
rect 378 267 384 268
rect 766 268 770 272
rect 774 268 778 272
rect 766 267 778 268
rect 159 263 160 267
rect 164 263 176 267
rect 180 263 312 267
rect 316 263 317 267
rect 159 262 317 263
rect 39 256 117 257
rect 39 252 40 256
rect 44 252 112 256
rect 116 252 117 256
rect 39 251 117 252
rect 271 239 309 240
rect 271 235 272 239
rect 276 235 304 239
rect 308 235 309 239
rect 271 234 309 235
rect -2 230 373 231
rect -2 226 0 230
rect 4 226 368 230
rect 372 226 373 230
rect -2 225 373 226
rect 47 177 149 178
rect 47 173 48 177
rect 52 173 144 177
rect 148 173 149 177
rect 47 172 149 173
rect 31 168 173 169
rect 31 164 32 168
rect 36 164 95 168
rect 100 164 168 168
rect 172 164 173 168
rect 31 163 173 164
rect 56 159 69 160
rect 56 155 57 159
rect 61 155 64 159
rect 68 155 69 159
rect 56 154 69 155
rect 159 157 317 158
rect 159 153 160 157
rect 164 153 176 157
rect 180 153 312 157
rect 316 153 317 157
rect 159 152 317 153
rect 39 146 117 147
rect 39 142 40 146
rect 44 142 112 146
rect 116 142 117 146
rect 39 141 117 142
rect 271 129 309 130
rect 271 125 272 129
rect 276 125 304 129
rect 308 125 309 129
rect 271 124 309 125
rect -2 120 373 121
rect -2 116 16 120
rect 20 116 368 120
rect 372 116 373 120
rect -2 115 373 116
rect 278 110 395 111
rect 278 106 279 110
rect 283 106 389 110
rect 393 106 395 110
rect 278 105 395 106
rect 79 101 384 102
rect 79 97 80 101
rect 84 97 379 101
rect 383 97 384 101
rect 79 96 384 97
rect 47 67 149 68
rect 47 63 48 67
rect 52 63 144 67
rect 148 63 149 67
rect 47 62 149 63
rect 378 62 384 63
rect 32 58 173 59
rect 32 54 33 58
rect 37 54 95 58
rect 100 54 168 58
rect 172 54 173 58
rect 32 53 173 54
rect 183 58 284 59
rect 183 56 279 58
rect 183 52 184 56
rect 188 54 279 56
rect 283 54 284 58
rect 378 58 379 62
rect 383 58 384 62
rect 378 57 384 58
rect 768 61 776 62
rect 768 57 769 61
rect 773 57 776 61
rect 188 53 284 54
rect 327 56 357 57
rect 768 56 774 57
rect 188 52 189 53
rect 183 51 189 52
rect 327 52 328 56
rect 332 52 352 56
rect 356 52 357 56
rect 327 51 357 52
rect 56 49 69 50
rect 56 45 57 49
rect 61 45 64 49
rect 68 45 69 49
rect 56 44 69 45
rect 159 47 317 48
rect 159 43 160 47
rect 164 43 176 47
rect 180 43 312 47
rect 316 43 317 47
rect 159 42 317 43
rect 39 36 117 37
rect 39 32 40 36
rect 44 32 112 36
rect 116 32 117 36
rect 39 31 117 32
rect 271 19 309 20
rect 271 15 272 19
rect 276 15 304 19
rect 308 15 309 19
rect 271 14 309 15
rect -2 10 373 11
rect -2 6 0 10
rect 4 6 368 10
rect 372 6 373 10
rect -2 5 373 6
use inv_1x  inv_1x_0
timestamp 1484418501
transform 1 0 265 0 1 884
box -6 -4 18 96
use yzdetect_8  yzdetect_8_0
timestamp 1484534894
transform 1 0 0 0 1 4
box -8 -4 28 756
use inv_1x_8  inv_1x_8_0
timestamp 1484534894
transform 1 0 32 0 1 4
box -6 -4 18 866
use inv_1x_8  inv_1x_8_1
timestamp 1484534894
transform 1 0 48 0 1 4
box -6 -4 18 866
use mux4_8_10space  mux4_8_10space_0
timestamp 1487099744
transform 1 0 58 0 1 0
box 0 0 112 870
use adder_8  adder_8_0
timestamp 1484427118
transform 1 0 168 0 1 4
box -6 -4 130 866
use mux3_1x_8  mux3_1x_8_0
timestamp 1484532969
transform 1 0 296 0 1 4
box -6 -4 82 976
use alu_ctl  alu_ctl_0
timestamp 1488311641
transform 1 0 378 0 1 0
box 0 0 400 980
<< labels >>
rlabel metal2 33 46 33 46 1 a0
rlabel metal2 49 46 49 46 1 b0
rlabel metal2 33 156 33 156 1 a1
rlabel metal2 49 156 49 156 1 b1
rlabel metal2 33 266 33 266 1 a2
rlabel metal2 49 266 49 266 1 b2
rlabel metal2 33 376 33 376 1 a3
rlabel metal2 49 376 49 376 1 b3
rlabel metal2 33 486 33 486 1 a4
rlabel metal2 49 486 49 486 1 b4
rlabel metal2 33 596 33 596 1 a5
rlabel metal3 -1 9 -1 9 1 result0
rlabel metal3 -1 119 -1 119 1 result1
rlabel metal3 -1 230 -1 230 1 result2
rlabel metal3 -1 340 -1 340 1 result3
rlabel metal3 -1 450 -1 450 1 result4
rlabel metal3 -1 560 -1 560 1 result5
rlabel metal3 -1 670 -1 670 1 result6
rlabel metal3 1 778 1 778 1 result7
rlabel m2contact 352 763 356 767 1 less
rlabel metal2 296 922 300 926 1 op0
rlabel metal2 328 922 332 926 1 op1
rlabel metal2 49 596 49 596 1 b5
rlabel metal2 33 706 33 706 1 a6
rlabel metal2 49 706 49 706 1 b6
rlabel metal2 33 816 33 816 1 a7
rlabel metal2 49 816 49 816 1 b7
rlabel metal2 9 370 9 370 1 zero
rlabel m3contact 161 44 161 44 1 muxy7
rlabel metal2 81 767 81 767 1 op6
rlabel metal2 89 767 89 767 1 op5
rlabel metal2 120 763 124 767 1 op4
rlabel metal2 136 763 140 767 1 op3
rlabel m3contact 98 56 98 56 1 mux4s1_0
rlabel metal2 146 61 146 61 1 mux4s0_0
rlabel m3contact 186 830 186 830 1 cout_adder_7
rlabel metal2 122 544 122 544 1 op4
rlabel metal2 90 325 90 325 1 op5
rlabel metal2 82 104 82 104 1 op6
rlabel metal2 281 106 281 106 1 op2
rlabel m2contact 554 45 554 45 1 Vdd!
rlabel m2contact 557 71 557 71 1 Gnd!
rlabel m3contact 771 699 771 699 1 funct_2
rlabel m3contact 771 489 771 489 1 funct_3
rlabel metal2 408 1 408 1 1 funct_0
rlabel metal2 719 1 719 1 1 alu_op_1
rlabel m3contact 772 269 772 269 1 funct_4
rlabel m3contact 773 920 773 920 1 funct_1
rlabel m3contact 381 470 381 470 1 alu_op_0
rlabel m3contact 771 59 771 59 1 funct_5
rlabel m3contact 186 53 186 53 1 op2
<< end >>
                                                                                                                                                                                                                                                                                                                                                                                                                                                alu_complete.mag                                                                                    0000644 �    Asz0000145 00000061004 13046424360 012136  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1486498032
<< nwell >>
rect 124 175 125 178
<< metal1 >>
rect 30 856 294 864
rect 348 803 352 807
rect -2 746 294 754
rect -2 662 366 664
rect -2 658 360 662
rect 364 658 366 662
rect -2 656 366 658
rect -2 636 294 644
rect -2 552 366 554
rect -2 548 360 552
rect 364 548 366 552
rect -2 546 366 548
rect -2 526 294 534
rect -2 442 366 444
rect -2 438 360 442
rect 364 438 366 442
rect -2 436 366 438
rect -2 416 294 424
rect -2 332 366 334
rect -2 328 360 332
rect 364 328 366 332
rect -2 326 366 328
rect -2 306 294 314
rect -2 222 366 224
rect -2 218 360 222
rect 364 218 366 222
rect -2 216 366 218
rect -2 196 294 204
rect -2 112 366 114
rect -2 108 360 112
rect 364 108 366 112
rect -2 106 366 108
rect -2 86 294 94
rect 356 33 363 37
rect -2 -4 294 4
<< m2contact >>
rect 344 803 348 807
rect 352 803 356 807
rect 360 768 364 772
rect 360 658 364 662
rect 360 548 364 552
rect 360 438 364 442
rect 360 328 364 332
rect 360 218 364 222
rect 360 108 364 112
rect 352 33 356 37
<< metal2 >>
rect 47 922 53 923
rect 47 918 48 922
rect 52 918 53 922
rect 47 917 53 918
rect 191 922 197 923
rect 191 918 192 922
rect 196 918 197 922
rect 288 918 292 922
rect 320 918 324 922
rect 191 917 197 918
rect 111 852 117 853
rect 111 848 112 852
rect 116 848 117 852
rect 111 847 117 848
rect 143 852 149 853
rect 143 848 144 852
rect 148 848 149 852
rect 143 847 149 848
rect 159 852 165 853
rect 159 848 160 852
rect 164 848 165 852
rect 159 847 165 848
rect 31 842 37 843
rect 31 838 32 842
rect 36 838 37 842
rect 31 837 37 838
rect 95 822 101 823
rect 95 818 96 822
rect 100 818 101 822
rect 95 817 101 818
rect 87 812 93 813
rect 87 808 88 812
rect 92 808 93 812
rect 96 809 100 817
rect 87 807 93 808
rect 112 801 116 847
rect 119 842 125 843
rect 119 838 120 842
rect 124 838 125 842
rect 119 837 125 838
rect 120 832 125 837
rect 144 818 148 847
rect 151 842 157 843
rect 151 838 152 842
rect 156 838 157 842
rect 151 837 157 838
rect 128 803 132 811
rect 127 802 133 803
rect 127 798 128 802
rect 132 798 133 802
rect 127 797 133 798
rect 152 793 156 837
rect 160 803 164 847
rect 167 812 173 813
rect 167 808 168 812
rect 172 808 173 812
rect 167 807 173 808
rect 15 782 21 783
rect 15 778 16 782
rect 20 778 21 782
rect 15 777 21 778
rect 0 673 4 706
rect 16 687 20 777
rect 111 742 117 743
rect 111 738 112 742
rect 116 738 117 742
rect 111 737 117 738
rect 143 742 149 743
rect 143 738 144 742
rect 148 738 149 742
rect 143 737 149 738
rect 159 742 165 743
rect 159 738 160 742
rect 164 738 165 742
rect 159 737 165 738
rect 31 732 37 733
rect 31 728 32 732
rect 36 728 37 732
rect 31 727 37 728
rect 95 712 101 713
rect 95 708 96 712
rect 100 708 101 712
rect 95 707 101 708
rect 87 702 93 703
rect 87 698 88 702
rect 92 698 93 702
rect 96 699 100 707
rect 87 697 93 698
rect 112 691 116 737
rect 119 732 125 733
rect 119 728 120 732
rect 124 728 125 732
rect 119 727 125 728
rect 120 722 125 727
rect 144 708 148 737
rect 151 732 157 733
rect 151 728 152 732
rect 156 728 157 732
rect 151 727 157 728
rect 128 693 132 701
rect 127 692 133 693
rect 127 688 128 692
rect 132 688 133 692
rect 127 687 133 688
rect 152 683 156 727
rect 160 693 164 737
rect 167 702 173 703
rect 167 698 168 702
rect 172 698 173 702
rect 167 697 173 698
rect -1 672 5 673
rect -1 668 0 672
rect 4 668 5 672
rect -1 667 5 668
rect 111 632 117 633
rect 111 628 112 632
rect 116 628 117 632
rect 111 627 117 628
rect 143 632 149 633
rect 143 628 144 632
rect 148 628 149 632
rect 143 627 149 628
rect 159 632 165 633
rect 159 628 160 632
rect 164 628 165 632
rect 159 627 165 628
rect 31 622 37 623
rect 31 618 32 622
rect 36 618 37 622
rect 31 617 37 618
rect 95 602 101 603
rect 95 598 96 602
rect 100 598 101 602
rect 95 597 101 598
rect 87 592 93 593
rect 87 588 88 592
rect 92 588 93 592
rect 96 589 100 597
rect 87 587 93 588
rect 112 581 116 627
rect 119 622 125 623
rect 119 618 120 622
rect 124 618 125 622
rect 119 617 125 618
rect 120 612 125 617
rect 144 598 148 627
rect 151 622 157 623
rect 151 618 152 622
rect 156 618 157 622
rect 151 617 157 618
rect 128 583 132 591
rect 127 582 133 583
rect 127 578 128 582
rect 132 578 133 582
rect 127 577 133 578
rect 152 573 156 617
rect 160 583 164 627
rect 167 592 173 593
rect 167 588 168 592
rect 172 588 173 592
rect 167 587 173 588
rect -1 562 5 563
rect -1 558 0 562
rect 4 558 5 562
rect -1 557 5 558
rect 0 484 4 557
rect 111 522 117 523
rect 111 518 112 522
rect 116 518 117 522
rect 111 517 117 518
rect 143 522 149 523
rect 143 518 144 522
rect 148 518 149 522
rect 143 517 149 518
rect 159 522 165 523
rect 159 518 160 522
rect 164 518 165 522
rect 159 517 165 518
rect 31 512 37 513
rect 31 508 32 512
rect 36 508 37 512
rect 31 507 37 508
rect 95 492 101 493
rect 95 488 96 492
rect 100 488 101 492
rect 95 487 101 488
rect 87 482 93 483
rect 87 478 88 482
rect 92 478 93 482
rect 96 479 100 487
rect 87 477 93 478
rect 112 471 116 517
rect 119 512 125 513
rect 119 508 120 512
rect 124 508 125 512
rect 119 507 125 508
rect 120 502 125 507
rect 144 488 148 517
rect 151 512 157 513
rect 151 508 152 512
rect 156 508 157 512
rect 151 507 157 508
rect 128 473 132 481
rect 127 472 133 473
rect 16 453 20 469
rect 127 468 128 472
rect 132 468 133 472
rect 127 467 133 468
rect 152 463 156 507
rect 160 473 164 517
rect 167 482 173 483
rect 167 478 168 482
rect 172 478 173 482
rect 167 477 173 478
rect 15 452 21 453
rect 15 448 16 452
rect 20 448 21 452
rect 15 447 21 448
rect 111 412 117 413
rect 111 408 112 412
rect 116 408 117 412
rect 111 407 117 408
rect 143 412 149 413
rect 143 408 144 412
rect 148 408 149 412
rect 143 407 149 408
rect 159 412 165 413
rect 159 408 160 412
rect 164 408 165 412
rect 159 407 165 408
rect 31 402 37 403
rect 31 398 32 402
rect 36 398 37 402
rect 31 397 37 398
rect 95 382 101 383
rect 95 378 96 382
rect 100 378 101 382
rect 95 377 101 378
rect 87 372 93 373
rect 87 368 88 372
rect 92 368 93 372
rect 96 369 100 377
rect 87 367 93 368
rect 8 363 12 367
rect 112 361 116 407
rect 119 402 125 403
rect 119 398 120 402
rect 124 398 125 402
rect 119 397 125 398
rect 120 392 125 397
rect 144 378 148 407
rect 151 402 157 403
rect 151 398 152 402
rect 156 398 157 402
rect 151 397 157 398
rect 128 363 132 371
rect 127 362 133 363
rect 127 358 128 362
rect 132 358 133 362
rect 127 357 133 358
rect 152 353 156 397
rect 160 363 164 407
rect 167 372 173 373
rect 167 368 168 372
rect 172 368 173 372
rect 167 367 173 368
rect 15 342 21 343
rect 15 338 16 342
rect 20 338 21 342
rect 15 337 21 338
rect 0 233 4 266
rect 16 247 20 337
rect 111 302 117 303
rect 111 298 112 302
rect 116 298 117 302
rect 111 297 117 298
rect 143 302 149 303
rect 143 298 144 302
rect 148 298 149 302
rect 143 297 149 298
rect 159 302 165 303
rect 159 298 160 302
rect 164 298 165 302
rect 159 297 165 298
rect 31 292 37 293
rect 31 288 32 292
rect 36 288 37 292
rect 95 272 101 273
rect 95 268 96 272
rect 100 268 101 272
rect 95 267 101 268
rect 87 262 93 263
rect 87 258 88 262
rect 92 258 93 262
rect 96 259 100 267
rect 87 257 93 258
rect 112 251 116 297
rect 119 292 125 293
rect 119 288 120 292
rect 124 288 125 292
rect 119 287 125 288
rect 120 285 125 287
rect 120 282 124 285
rect 144 268 148 297
rect 151 292 157 293
rect 151 288 152 292
rect 156 288 157 292
rect 151 287 157 288
rect 128 253 132 261
rect 127 252 133 253
rect 127 248 128 252
rect 132 248 133 252
rect 127 247 133 248
rect 152 243 156 287
rect 160 253 164 297
rect 167 262 173 263
rect 167 258 168 262
rect 172 258 173 262
rect 167 257 173 258
rect -1 232 5 233
rect -1 228 0 232
rect 4 228 5 232
rect -1 227 5 228
rect 111 192 117 193
rect 111 188 112 192
rect 116 188 117 192
rect 111 187 117 188
rect 143 192 149 193
rect 143 188 144 192
rect 148 188 149 192
rect 143 187 149 188
rect 159 192 165 193
rect 159 188 160 192
rect 164 188 165 192
rect 159 187 165 188
rect 95 162 101 163
rect 95 158 96 162
rect 100 158 101 162
rect 95 157 101 158
rect 87 152 93 153
rect 87 148 88 152
rect 92 148 93 152
rect 96 149 100 157
rect 87 147 93 148
rect 112 141 116 187
rect 119 182 125 183
rect 119 178 120 182
rect 124 178 125 182
rect 119 177 125 178
rect 120 175 125 177
rect 120 172 124 175
rect 144 158 148 187
rect 151 182 157 183
rect 151 178 152 182
rect 156 178 157 182
rect 151 177 157 178
rect 128 143 132 151
rect 127 142 133 143
rect 127 138 128 142
rect 132 138 133 142
rect 127 137 133 138
rect 152 133 156 177
rect 160 143 164 187
rect 167 152 173 153
rect 167 148 168 152
rect 172 148 173 152
rect 167 147 173 148
rect 15 122 21 123
rect 15 118 16 122
rect 20 118 21 122
rect 15 117 21 118
rect 0 13 4 46
rect 16 27 20 117
rect 111 82 117 83
rect 111 78 112 82
rect 116 78 117 82
rect 111 77 117 78
rect 143 82 149 83
rect 143 78 144 82
rect 148 78 149 82
rect 143 77 149 78
rect 159 82 165 83
rect 159 78 160 82
rect 164 78 165 82
rect 159 77 165 78
rect 31 72 37 73
rect 31 68 32 72
rect 36 68 37 72
rect 31 67 37 68
rect 95 52 101 53
rect 95 48 96 52
rect 100 48 101 52
rect 95 47 101 48
rect 87 42 93 43
rect 87 38 88 42
rect 92 38 93 42
rect 96 39 100 47
rect 87 37 93 38
rect 112 31 116 77
rect 119 72 125 73
rect 119 68 120 72
rect 124 68 125 72
rect 119 67 125 68
rect 120 65 125 67
rect 120 62 124 65
rect 144 48 148 77
rect 151 72 157 73
rect 151 68 152 72
rect 156 68 157 72
rect 151 67 157 68
rect 128 33 132 41
rect 127 32 133 33
rect 127 28 128 32
rect 132 28 133 32
rect 127 27 133 28
rect 152 23 156 67
rect 160 33 164 77
rect 167 42 173 43
rect 167 38 168 42
rect 172 38 173 42
rect 167 37 173 38
rect 176 23 180 50
rect 192 23 196 917
rect 263 852 269 853
rect 263 848 264 852
rect 268 848 269 852
rect 263 847 269 848
rect 343 852 349 853
rect 343 848 344 852
rect 348 848 349 852
rect 343 847 349 848
rect 264 782 268 847
rect 303 822 309 823
rect 303 818 304 822
rect 308 818 309 822
rect 303 817 309 818
rect 304 805 308 817
rect 344 807 348 847
rect 312 803 316 807
rect 311 802 317 803
rect 311 798 312 802
rect 316 798 317 802
rect 311 797 317 798
rect 263 742 269 743
rect 263 738 264 742
rect 268 738 269 742
rect 263 737 269 738
rect 343 742 349 743
rect 343 738 344 742
rect 348 738 349 742
rect 343 737 349 738
rect 264 672 268 737
rect 303 712 309 713
rect 303 708 304 712
rect 308 708 309 712
rect 344 710 348 737
rect 303 707 309 708
rect 304 695 308 707
rect 312 693 316 697
rect 311 692 317 693
rect 311 688 312 692
rect 316 688 317 692
rect 311 687 317 688
rect 263 632 269 633
rect 263 628 264 632
rect 268 628 269 632
rect 263 627 269 628
rect 343 632 349 633
rect 343 628 344 632
rect 348 628 349 632
rect 343 627 349 628
rect 264 562 268 627
rect 303 602 309 603
rect 303 598 304 602
rect 308 598 309 602
rect 344 600 348 627
rect 303 597 309 598
rect 304 585 308 597
rect 312 583 316 587
rect 311 582 317 583
rect 311 578 312 582
rect 316 578 317 582
rect 311 577 317 578
rect 263 522 269 523
rect 263 518 264 522
rect 268 518 269 522
rect 263 517 269 518
rect 343 522 349 523
rect 343 518 344 522
rect 348 518 349 522
rect 343 517 349 518
rect 264 452 268 517
rect 303 492 309 493
rect 303 488 304 492
rect 308 488 309 492
rect 344 490 348 517
rect 303 487 309 488
rect 304 475 308 487
rect 312 473 316 477
rect 311 472 317 473
rect 311 468 312 472
rect 316 468 317 472
rect 311 467 317 468
rect 263 412 269 413
rect 263 408 264 412
rect 268 408 269 412
rect 263 407 269 408
rect 343 412 349 413
rect 343 408 344 412
rect 348 408 349 412
rect 343 407 349 408
rect 264 342 268 407
rect 303 382 309 383
rect 303 378 304 382
rect 308 378 309 382
rect 344 380 348 407
rect 303 377 309 378
rect 304 365 308 377
rect 312 363 316 367
rect 311 362 317 363
rect 311 358 312 362
rect 316 358 317 362
rect 311 357 317 358
rect 263 302 269 303
rect 263 298 264 302
rect 268 298 269 302
rect 263 297 269 298
rect 343 302 349 303
rect 343 298 344 302
rect 348 298 349 302
rect 343 297 349 298
rect 264 232 268 297
rect 303 272 309 273
rect 303 268 304 272
rect 308 268 309 272
rect 344 270 348 297
rect 303 267 309 268
rect 304 255 308 267
rect 312 253 316 257
rect 311 252 317 253
rect 311 248 312 252
rect 316 248 317 252
rect 311 247 317 248
rect 263 192 269 193
rect 263 188 264 192
rect 268 188 269 192
rect 263 187 269 188
rect 343 192 349 193
rect 343 188 344 192
rect 348 188 349 192
rect 343 187 349 188
rect 264 122 268 187
rect 303 162 309 163
rect 303 158 304 162
rect 308 158 309 162
rect 344 160 348 187
rect 303 157 309 158
rect 304 145 308 157
rect 312 143 316 147
rect 311 142 317 143
rect 311 138 312 142
rect 316 138 317 142
rect 311 137 317 138
rect 263 82 269 83
rect 263 78 264 82
rect 268 78 269 82
rect 263 77 269 78
rect 343 82 349 83
rect 343 78 344 82
rect 348 78 349 82
rect 343 77 349 78
rect 175 22 181 23
rect 175 18 176 22
rect 180 18 181 22
rect 175 17 181 18
rect 191 22 197 23
rect 191 18 192 22
rect 196 18 197 22
rect 191 17 197 18
rect -1 12 5 13
rect 264 12 268 77
rect 303 52 309 53
rect 303 48 304 52
rect 308 48 309 52
rect 344 50 348 77
rect 303 47 309 48
rect 304 35 308 47
rect 352 37 356 803
rect 360 772 364 806
rect 384 783 388 810
rect 383 782 389 783
rect 383 778 384 782
rect 388 778 389 782
rect 383 777 389 778
rect 360 662 364 696
rect 384 673 388 700
rect 383 672 389 673
rect 383 668 384 672
rect 388 668 389 672
rect 383 667 389 668
rect 360 552 364 586
rect 384 563 388 590
rect 383 562 389 563
rect 383 558 384 562
rect 388 558 389 562
rect 383 557 389 558
rect 360 442 364 476
rect 384 453 388 480
rect 383 452 389 453
rect 383 448 384 452
rect 388 448 389 452
rect 383 447 389 448
rect 360 332 364 366
rect 384 343 388 370
rect 383 342 389 343
rect 383 338 384 342
rect 388 338 389 342
rect 383 337 389 338
rect 360 222 364 256
rect 384 233 388 260
rect 383 232 389 233
rect 383 228 384 232
rect 388 228 389 232
rect 383 227 389 228
rect 360 112 364 146
rect 384 123 388 150
rect 383 122 389 123
rect 383 118 384 122
rect 388 118 389 122
rect 383 117 389 118
rect 312 33 316 37
rect 311 32 317 33
rect 311 28 312 32
rect 316 28 317 32
rect 311 27 317 28
rect 384 13 388 40
rect 383 12 389 13
rect -1 8 0 12
rect 4 8 5 12
rect -1 7 5 8
rect 383 8 384 12
rect 388 8 389 12
rect 383 7 389 8
<< m3contact >>
rect 48 918 52 922
rect 192 918 196 922
rect 112 848 116 852
rect 144 848 148 852
rect 160 848 164 852
rect 32 838 36 842
rect 96 818 100 822
rect 88 808 92 812
rect 120 838 124 842
rect 152 838 156 842
rect 128 798 132 802
rect 168 808 172 812
rect 16 778 20 782
rect 112 738 116 742
rect 144 738 148 742
rect 160 738 164 742
rect 32 728 36 732
rect 96 708 100 712
rect 88 698 92 702
rect 120 728 124 732
rect 152 728 156 732
rect 128 688 132 692
rect 168 698 172 702
rect 0 668 4 672
rect 112 628 116 632
rect 144 628 148 632
rect 160 628 164 632
rect 32 618 36 622
rect 96 598 100 602
rect 88 588 92 592
rect 120 618 124 622
rect 152 618 156 622
rect 128 578 132 582
rect 168 588 172 592
rect 0 558 4 562
rect 112 518 116 522
rect 144 518 148 522
rect 160 518 164 522
rect 32 508 36 512
rect 96 488 100 492
rect 88 478 92 482
rect 120 508 124 512
rect 152 508 156 512
rect 128 468 132 472
rect 168 478 172 482
rect 16 448 20 452
rect 112 408 116 412
rect 144 408 148 412
rect 160 408 164 412
rect 32 398 36 402
rect 96 378 100 382
rect 88 368 92 372
rect 120 398 124 402
rect 152 398 156 402
rect 128 358 132 362
rect 168 368 172 372
rect 16 338 20 342
rect 112 298 116 302
rect 144 298 148 302
rect 160 298 164 302
rect 32 288 36 292
rect 96 268 100 272
rect 88 258 92 262
rect 120 288 124 292
rect 152 288 156 292
rect 128 248 132 252
rect 168 258 172 262
rect 0 228 4 232
rect 112 188 116 192
rect 144 188 148 192
rect 160 188 164 192
rect 96 158 100 162
rect 88 148 92 152
rect 120 178 124 182
rect 152 178 156 182
rect 128 138 132 142
rect 168 148 172 152
rect 16 118 20 122
rect 112 78 116 82
rect 144 78 148 82
rect 160 78 164 82
rect 32 68 36 72
rect 96 48 100 52
rect 88 38 92 42
rect 120 68 124 72
rect 152 68 156 72
rect 128 28 132 32
rect 168 38 172 42
rect 264 848 268 852
rect 344 848 348 852
rect 304 818 308 822
rect 312 798 316 802
rect 264 738 268 742
rect 344 738 348 742
rect 304 708 308 712
rect 312 688 316 692
rect 264 628 268 632
rect 344 628 348 632
rect 304 598 308 602
rect 312 578 316 582
rect 264 518 268 522
rect 344 518 348 522
rect 304 488 308 492
rect 312 468 316 472
rect 264 408 268 412
rect 344 408 348 412
rect 304 378 308 382
rect 312 358 316 362
rect 264 298 268 302
rect 344 298 348 302
rect 304 268 308 272
rect 312 248 316 252
rect 264 188 268 192
rect 344 188 348 192
rect 304 158 308 162
rect 312 138 316 142
rect 264 78 268 82
rect 344 78 348 82
rect 176 18 180 22
rect 192 18 196 22
rect 304 48 308 52
rect 384 778 388 782
rect 384 668 388 672
rect 384 558 388 562
rect 384 448 388 452
rect 384 338 388 342
rect 384 228 388 232
rect 384 118 388 122
rect 312 28 316 32
rect 0 8 4 12
rect 384 8 388 12
<< metal3 >>
rect 47 922 197 923
rect 47 918 48 922
rect 52 918 192 922
rect 196 918 197 922
rect 47 917 197 918
rect -17 852 165 853
rect -17 848 112 852
rect 116 848 144 852
rect 148 848 160 852
rect 164 848 165 852
rect -17 847 165 848
rect 263 852 349 853
rect 263 848 264 852
rect 268 848 344 852
rect 348 848 349 852
rect 263 847 349 848
rect -17 842 157 843
rect -17 838 32 842
rect 36 838 120 842
rect 124 838 152 842
rect 156 838 157 842
rect -17 837 157 838
rect 95 822 309 823
rect 95 818 96 822
rect 100 818 304 822
rect 308 818 309 822
rect 95 817 309 818
rect 87 812 173 813
rect 87 808 88 812
rect 92 808 168 812
rect 172 808 173 812
rect 87 807 173 808
rect 127 802 317 803
rect 127 798 128 802
rect 132 798 312 802
rect 316 798 317 802
rect 127 797 317 798
rect -17 782 389 783
rect -17 778 16 782
rect 20 778 384 782
rect 388 778 389 782
rect -17 777 389 778
rect -17 742 165 743
rect -17 738 112 742
rect 116 738 144 742
rect 148 738 160 742
rect 164 738 165 742
rect -17 737 165 738
rect 263 742 349 743
rect 263 738 264 742
rect 268 738 344 742
rect 348 738 349 742
rect 263 737 349 738
rect -17 732 157 733
rect -17 728 32 732
rect 36 728 120 732
rect 124 728 152 732
rect 156 728 157 732
rect -17 727 157 728
rect 95 712 309 713
rect 95 708 96 712
rect 100 708 304 712
rect 308 708 309 712
rect 95 707 309 708
rect 87 702 173 703
rect 87 698 88 702
rect 92 698 168 702
rect 172 698 173 702
rect 87 697 173 698
rect 127 692 317 693
rect 127 688 128 692
rect 132 688 312 692
rect 316 688 317 692
rect 127 687 317 688
rect -17 672 389 673
rect -17 668 0 672
rect 4 668 384 672
rect 388 668 389 672
rect -17 667 389 668
rect -17 632 165 633
rect -17 628 112 632
rect 116 628 144 632
rect 148 628 160 632
rect 164 628 165 632
rect -17 627 165 628
rect 263 632 349 633
rect 263 628 264 632
rect 268 628 344 632
rect 348 628 349 632
rect 263 627 349 628
rect -17 622 157 623
rect -17 618 32 622
rect 36 618 120 622
rect 124 618 152 622
rect 156 618 157 622
rect -17 617 157 618
rect 95 602 309 603
rect 95 598 96 602
rect 100 598 304 602
rect 308 598 309 602
rect 95 597 309 598
rect 87 592 173 593
rect 87 588 88 592
rect 92 588 168 592
rect 172 588 173 592
rect 87 587 173 588
rect 127 582 317 583
rect 127 578 128 582
rect 132 578 312 582
rect 316 578 317 582
rect 127 577 317 578
rect -17 562 389 563
rect -17 558 0 562
rect 4 558 384 562
rect 388 558 389 562
rect -17 557 389 558
rect -17 522 165 523
rect -17 518 112 522
rect 116 518 144 522
rect 148 518 160 522
rect 164 518 165 522
rect -17 517 165 518
rect 263 522 349 523
rect 263 518 264 522
rect 268 518 344 522
rect 348 518 349 522
rect 263 517 349 518
rect -17 512 157 513
rect -17 508 32 512
rect 36 508 120 512
rect 124 508 152 512
rect 156 508 157 512
rect -17 507 157 508
rect 95 492 309 493
rect 95 488 96 492
rect 100 488 304 492
rect 308 488 309 492
rect 95 487 309 488
rect 87 482 173 483
rect 87 478 88 482
rect 92 478 168 482
rect 172 478 173 482
rect 87 477 173 478
rect 127 472 317 473
rect 127 468 128 472
rect 132 468 312 472
rect 316 468 317 472
rect 127 467 317 468
rect -17 452 389 453
rect -17 448 16 452
rect 20 448 384 452
rect 388 448 389 452
rect -17 447 389 448
rect -17 412 165 413
rect -17 408 112 412
rect 116 408 144 412
rect 148 408 160 412
rect 164 408 165 412
rect -17 407 165 408
rect 263 412 349 413
rect 263 408 264 412
rect 268 408 344 412
rect 348 408 349 412
rect 263 407 349 408
rect -17 402 157 403
rect -17 398 32 402
rect 36 398 120 402
rect 124 398 152 402
rect 156 398 157 402
rect -17 397 157 398
rect 95 382 309 383
rect 95 378 96 382
rect 100 378 304 382
rect 308 378 309 382
rect 95 377 309 378
rect 87 372 173 373
rect 87 368 88 372
rect 92 368 168 372
rect 172 368 173 372
rect 87 367 173 368
rect 127 362 317 363
rect 127 358 128 362
rect 132 358 312 362
rect 316 358 317 362
rect 127 357 317 358
rect -17 342 389 343
rect -17 338 16 342
rect 20 338 384 342
rect 388 338 389 342
rect -17 337 389 338
rect -17 302 165 303
rect -17 298 112 302
rect 116 298 144 302
rect 148 298 160 302
rect 164 298 165 302
rect -17 297 165 298
rect 263 302 349 303
rect 263 298 264 302
rect 268 298 344 302
rect 348 298 349 302
rect 263 297 349 298
rect -17 292 157 293
rect -17 288 32 292
rect 36 288 120 292
rect 124 288 152 292
rect 156 288 157 292
rect -17 287 21 288
rect 85 287 157 288
rect 95 272 309 273
rect 95 268 96 272
rect 100 268 304 272
rect 308 268 309 272
rect 95 267 309 268
rect 87 262 173 263
rect 87 258 88 262
rect 92 258 168 262
rect 172 258 173 262
rect 87 257 173 258
rect 127 252 317 253
rect 127 248 128 252
rect 132 248 312 252
rect 316 248 317 252
rect 127 247 317 248
rect -17 232 389 233
rect -17 228 0 232
rect 4 228 384 232
rect 388 228 389 232
rect -17 227 389 228
rect -17 192 165 193
rect -17 188 112 192
rect 116 188 144 192
rect 148 188 160 192
rect 164 188 165 192
rect -17 187 165 188
rect 263 192 349 193
rect 263 188 264 192
rect 268 188 344 192
rect 348 188 349 192
rect 263 187 349 188
rect -17 182 157 183
rect -17 178 120 182
rect 124 178 152 182
rect 156 178 157 182
rect -17 177 157 178
rect 95 162 309 163
rect 95 158 96 162
rect 100 158 304 162
rect 308 158 309 162
rect 95 157 309 158
rect 87 152 173 153
rect 87 148 88 152
rect 92 148 168 152
rect 172 148 173 152
rect 87 147 173 148
rect 127 142 317 143
rect 127 138 128 142
rect 132 138 312 142
rect 316 138 317 142
rect 127 137 317 138
rect -17 122 389 123
rect -17 118 16 122
rect 20 118 384 122
rect 388 118 389 122
rect -17 117 389 118
rect -17 82 165 83
rect -17 78 112 82
rect 116 78 144 82
rect 148 78 160 82
rect 164 78 165 82
rect -17 77 165 78
rect 263 82 349 83
rect 263 78 264 82
rect 268 78 344 82
rect 348 78 349 82
rect 263 77 349 78
rect -17 72 157 73
rect -17 68 32 72
rect 36 68 120 72
rect 124 68 152 72
rect 156 68 157 72
rect -17 67 157 68
rect 95 52 309 53
rect 95 48 96 52
rect 100 48 304 52
rect 308 48 309 52
rect 95 47 309 48
rect 87 42 173 43
rect 87 38 88 42
rect 92 38 168 42
rect 172 38 173 42
rect 87 37 173 38
rect 127 32 317 33
rect 127 28 128 32
rect 132 28 312 32
rect 316 28 317 32
rect 127 27 317 28
rect 175 22 197 23
rect 175 18 176 22
rect 180 18 192 22
rect 196 18 197 22
rect 175 17 197 18
rect -17 12 389 13
rect -17 8 0 12
rect 4 8 384 12
rect 388 8 389 12
rect -17 7 389 8
use yzdetect_8  yzdetect_8_0
timestamp 1484534894
transform 1 0 0 0 1 0
box -8 -4 28 756
use condinv  condinv_0
timestamp 1484534894
transform 1 0 32 0 1 0
box -6 -4 66 976
use and2_1x_8  and2_1x_8_0
timestamp 1486497882
transform 1 0 90 0 1 -4
box 0 0 40 870
use or2_1x_8  or2_1x_8_0
timestamp 1484433330
transform 1 0 128 0 1 0
box -6 -4 34 866
use adder_8  adder_8_0
timestamp 1484427118
transform 1 0 160 0 1 0
box -6 -4 130 866
use mux4_1x_8  mux4_1x_8_0
timestamp 1484532969
transform 1 0 288 0 1 0
box -6 -4 106 976
<< labels >>
rlabel metal3 -15 10 -15 10 3 result_0_
rlabel metal3 -15 69 -15 69 3 b_0_
rlabel metal3 -14 80 -14 80 3 a_0_
rlabel metal3 -14 120 -14 120 3 result_1_
rlabel metal3 -14 180 -14 180 3 b_1_
rlabel metal3 -14 190 -14 190 3 a_1_
rlabel metal3 -14 230 -14 230 3 result_2_
rlabel metal3 -14 290 -14 290 3 b_2_
rlabel metal3 -13 300 -13 300 3 a_2_
rlabel metal3 -13 399 -13 399 3 b_3_
rlabel metal3 -15 510 -15 510 3 b_4_
rlabel metal3 -14 520 -14 520 3 a_4_
rlabel metal3 -14 560 -14 560 3 result_5_
rlabel metal3 -13 620 -13 620 3 b_5_
rlabel metal3 -14 630 -14 630 3 a_5_
rlabel metal3 -14 669 -14 669 3 result_6_
rlabel metal3 -13 730 -13 730 3 b_6_
rlabel metal3 -13 739 -13 739 3 a_6_
rlabel metal3 -14 780 -14 780 3 result_7_
rlabel metal3 -14 839 -14 839 3 b_7_
rlabel metal3 -14 850 -14 850 3 a_7_
rlabel metal3 55 920 55 920 1 alucontrol_2_
rlabel metal1 33 860 33 860 1 Vdd!
rlabel metal1 6 549 6 549 1 Gnd!
rlabel metal1 6 530 6 530 1 Vdd!
rlabel metal1 4 219 4 219 1 Gnd!
rlabel metal1 2 200 2 200 1 Vdd!
rlabel metal1 3 109 3 109 1 Gnd!
rlabel metal1 1 90 1 90 1 Vdd!
rlabel metal1 3 -1 3 -1 1 Gnd!
rlabel metal2 288 918 292 922 1 alucontrol_0_
rlabel metal2 320 918 324 922 1 alucontrol_1_
rlabel metal1 3 310 3 310 1 Vdd!
rlabel metal1 5 330 5 330 1 Gnd!
rlabel metal1 4 419 4 419 1 Vdd!
rlabel metal1 5 440 5 440 1 Gnd!
rlabel metal1 2 640 2 640 1 Vdd!
rlabel metal1 1 659 1 659 1 Gnd!
rlabel metal1 2 749 2 749 1 Vdd!
rlabel metal2 8 363 12 367 1 zero
rlabel metal3 -13 340 -13 340 3 result_3_
rlabel metal3 -14 450 -14 450 3 result_4_
rlabel metal3 -14 410 -14 410 3 a_3_
<< end >>
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            alu_ctl.mag                                                                                         0000644 �    Asz0000145 00000112363 13055352531 011115  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1488311641
<< metal1 >>
rect 30 925 370 940
rect 55 900 345 915
rect 55 887 345 893
rect 202 868 269 871
rect 162 841 177 844
rect 107 798 117 801
rect 195 798 237 801
rect 30 787 370 793
rect 147 741 157 744
rect 90 721 129 724
rect 217 723 222 732
rect 55 687 345 693
rect 130 648 134 657
rect 195 651 205 654
rect 218 651 222 654
rect 218 648 229 651
rect 266 648 279 653
rect 291 651 317 654
rect 210 638 229 641
rect 106 628 113 636
rect 266 631 273 636
rect 234 628 273 631
rect 30 587 370 593
rect 106 578 117 581
rect 186 548 197 551
rect 234 528 277 531
rect 290 528 294 537
rect 129 519 134 523
rect 211 519 221 522
rect 55 487 345 493
rect 90 478 101 481
rect 107 451 125 454
rect 250 451 277 454
rect 162 450 197 451
rect 162 448 221 450
rect 194 447 221 448
rect 202 438 213 441
rect 295 431 302 436
rect 218 428 229 431
rect 295 428 309 431
rect 235 398 261 401
rect 30 387 370 393
rect 255 344 262 352
rect 98 338 109 341
rect 218 321 241 324
rect 258 312 262 327
rect 120 298 133 301
rect 55 287 345 293
rect 154 278 164 282
rect 106 248 149 251
rect 247 231 254 236
rect 247 228 269 231
rect 30 187 370 193
rect 186 178 195 182
rect 98 145 113 148
rect 306 128 310 137
rect 234 121 269 122
rect 219 119 269 121
rect 219 118 237 119
rect 55 87 345 93
rect 55 65 345 80
rect 30 40 370 55
<< metal2 >>
rect 18 977 45 980
rect 314 977 357 980
rect 18 868 21 977
rect 18 3 21 261
rect 30 40 45 940
rect 55 65 70 915
rect 106 861 109 921
rect 194 868 205 871
rect 98 858 109 861
rect 98 851 101 858
rect 90 498 93 721
rect 98 311 101 801
rect 106 678 109 858
rect 226 851 277 854
rect 138 731 141 851
rect 130 728 141 731
rect 98 308 109 311
rect 98 251 101 261
rect 106 231 109 308
rect 98 228 109 231
rect 114 228 117 691
rect 130 578 133 651
rect 138 521 141 728
rect 138 518 149 521
rect 130 508 141 511
rect 122 368 125 501
rect 122 341 125 351
rect 130 341 133 508
rect 146 471 149 518
rect 122 338 133 341
rect 138 468 149 471
rect 122 258 125 338
rect 98 145 101 228
rect 106 158 109 201
rect 122 135 125 151
rect 130 125 133 301
rect 138 248 141 468
rect 154 278 157 744
rect 162 478 165 844
rect 162 331 165 451
rect 170 348 173 531
rect 178 378 181 721
rect 202 651 205 724
rect 210 688 213 732
rect 226 718 229 851
rect 186 548 189 651
rect 202 588 205 631
rect 162 328 173 331
rect 146 248 165 251
rect 162 241 165 248
rect 170 245 173 328
rect 178 278 181 371
rect 162 238 181 241
rect 186 178 189 341
rect 178 115 181 161
rect 194 148 197 501
rect 210 391 213 661
rect 218 428 221 701
rect 234 628 237 801
rect 250 698 253 725
rect 202 388 213 391
rect 202 278 205 388
rect 218 321 221 331
rect 226 318 229 591
rect 266 488 269 651
rect 250 441 253 454
rect 274 451 277 701
rect 282 647 285 661
rect 290 491 293 531
rect 298 528 301 921
rect 314 728 317 977
rect 306 688 309 701
rect 314 698 317 722
rect 290 488 301 491
rect 274 448 285 451
rect 242 438 253 441
rect 242 338 245 438
rect 258 348 261 431
rect 202 228 205 241
rect 210 115 213 291
rect 226 238 229 281
rect 234 231 237 251
rect 218 228 237 231
rect 242 228 245 261
rect 274 253 278 262
rect 290 228 293 401
rect 218 141 221 228
rect 298 171 301 488
rect 314 378 317 654
rect 306 178 309 261
rect 298 168 309 171
rect 218 138 229 141
rect 274 118 277 131
rect 106 58 109 101
rect 282 58 285 151
rect 306 128 309 168
rect 314 3 317 241
rect 330 65 345 915
rect 355 40 370 940
rect 18 0 45 3
rect 314 0 357 3
<< metal3 >>
rect 0 917 110 922
rect 297 917 400 922
rect 17 867 198 872
rect 137 847 182 852
rect 97 797 118 802
rect 217 727 318 732
rect 177 717 230 722
rect 0 697 150 702
rect 217 697 400 702
rect 113 687 310 692
rect 201 663 206 672
rect 201 662 214 663
rect 201 657 286 662
rect 185 647 230 652
rect 121 637 230 642
rect 105 627 238 632
rect 201 587 302 592
rect 105 577 134 582
rect 169 527 238 532
rect 129 517 222 522
rect 89 497 126 502
rect 0 487 270 492
rect 297 487 400 492
rect 89 477 166 482
rect 0 467 142 472
rect 201 437 246 442
rect 257 427 310 432
rect 121 367 182 372
rect 105 332 110 342
rect 121 337 246 342
rect 105 327 222 332
rect 89 317 230 322
rect 257 317 310 322
rect 209 287 270 292
rect 177 277 230 282
rect 265 272 270 287
rect 0 267 254 272
rect 265 267 400 272
rect 17 257 126 262
rect 217 257 310 262
rect 137 247 238 252
rect 201 237 318 242
rect 161 227 246 232
rect 265 227 286 232
rect 105 157 182 162
rect 121 147 198 152
rect 193 127 278 132
rect 273 117 294 122
rect 0 57 110 62
rect 281 57 400 62
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_0
timestamp 1488311641
transform 1 0 37 0 1 932
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_1
timestamp 1488311641
transform 1 0 362 0 1 932
box -7 -7 7 7
use $$M3_M2  $$M3_M2_0
timestamp 1488311641
transform 1 0 108 0 1 920
box -3 -3 3 3
use $$M3_M2  $$M3_M2_1
timestamp 1488311641
transform 1 0 300 0 1 920
box -3 -3 3 3
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_2
timestamp 1488311641
transform 1 0 62 0 1 907
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_3
timestamp 1488311641
transform 1 0 337 0 1 907
box -7 -7 7 7
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_0
timestamp 1488311641
transform 1 0 62 0 1 890
box -7 -2 7 2
use $$M3_M2  $$M3_M2_2
timestamp 1488311641
transform 1 0 20 0 1 870
box -3 -3 3 3
use $$M2_M1  $$M2_M1_0
timestamp 1488311641
transform 1 0 100 0 1 853
box -2 -2 2 2
use $$M3_M2  $$M3_M2_3
timestamp 1488311641
transform 1 0 100 0 1 800
box -3 -3 3 3
use $$M2_M1  $$M2_M1_1
timestamp 1488311641
transform 1 0 116 0 1 800
box -2 -2 2 2
use $$M3_M2  $$M3_M2_4
timestamp 1488311641
transform 1 0 116 0 1 800
box -3 -3 3 3
use $$M3_M2  $$M3_M2_5
timestamp 1488311641
transform 1 0 140 0 1 850
box -3 -3 3 3
use $$M2_M1  $$M2_M1_2
timestamp 1488311641
transform 1 0 164 0 1 843
box -2 -2 2 2
use $$M2_M1  $$M2_M1_3
timestamp 1488311641
transform 1 0 196 0 1 869
box -2 -2 2 2
use $$M3_M2  $$M3_M2_6
timestamp 1488311641
transform 1 0 196 0 1 870
box -3 -3 3 3
use $$M2_M1  $$M2_M1_4
timestamp 1488311641
transform 1 0 204 0 1 870
box -2 -2 2 2
use $$M2_M1  $$M2_M1_5
timestamp 1488311641
transform 1 0 180 0 1 852
box -2 -2 2 2
use $$M3_M2  $$M3_M2_7
timestamp 1488311641
transform 1 0 180 0 1 850
box -3 -3 3 3
use $$M2_M1  $$M2_M1_6
timestamp 1488311641
transform 1 0 236 0 1 800
box -2 -2 2 2
use $$M2_M1  $$M2_M1_7
timestamp 1488311641
transform 1 0 276 0 1 853
box -2 -2 2 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_1
timestamp 1488311641
transform 1 0 337 0 1 890
box -7 -2 7 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_2
timestamp 1488311641
transform 1 0 37 0 1 790
box -7 -2 7 2
use FILL  FILL_0
timestamp 1488311641
transform 1 0 80 0 -1 890
box -8 -3 16 105
use FILL  FILL_1
timestamp 1488311641
transform 1 0 88 0 -1 890
box -8 -3 16 105
use INVX2  INVX2_0
timestamp 1488311641
transform 1 0 96 0 -1 890
box -9 -3 26 105
use FILL  FILL_2
timestamp 1488311641
transform 1 0 112 0 -1 890
box -8 -3 16 105
use FILL  FILL_3
timestamp 1488311641
transform 1 0 120 0 -1 890
box -8 -3 16 105
use FILL  FILL_4
timestamp 1488311641
transform 1 0 128 0 -1 890
box -8 -3 16 105
use FILL  FILL_5
timestamp 1488311641
transform 1 0 136 0 -1 890
box -8 -3 16 105
use FILL  FILL_6
timestamp 1488311641
transform 1 0 144 0 -1 890
box -8 -3 16 105
use FILL  FILL_7
timestamp 1488311641
transform 1 0 152 0 -1 890
box -8 -3 16 105
use FILL  FILL_8
timestamp 1488311641
transform 1 0 160 0 -1 890
box -8 -3 16 105
use AOI21X1  AOI21X1_0
timestamp 1488311641
transform 1 0 168 0 -1 890
box -7 -3 39 105
use FILL  FILL_9
timestamp 1488311641
transform 1 0 200 0 -1 890
box -8 -3 16 105
use FILL  FILL_10
timestamp 1488311641
transform 1 0 208 0 -1 890
box -8 -3 16 105
use FILL  FILL_11
timestamp 1488311641
transform 1 0 216 0 -1 890
box -8 -3 16 105
use FILL  FILL_12
timestamp 1488311641
transform 1 0 224 0 -1 890
box -8 -3 16 105
use FILL  FILL_13
timestamp 1488311641
transform 1 0 232 0 -1 890
box -8 -3 16 105
use FILL  FILL_14
timestamp 1488311641
transform 1 0 240 0 -1 890
box -8 -3 16 105
use FILL  FILL_15
timestamp 1488311641
transform 1 0 248 0 -1 890
box -8 -3 16 105
use FILL  FILL_16
timestamp 1488311641
transform 1 0 256 0 -1 890
box -8 -3 16 105
use INVX2  INVX2_1
timestamp 1488311641
transform -1 0 280 0 -1 890
box -9 -3 26 105
use FILL  FILL_17
timestamp 1488311641
transform 1 0 280 0 -1 890
box -8 -3 16 105
use FILL  FILL_18
timestamp 1488311641
transform 1 0 288 0 -1 890
box -8 -3 16 105
use FILL  FILL_19
timestamp 1488311641
transform 1 0 296 0 -1 890
box -8 -3 16 105
use FILL  FILL_20
timestamp 1488311641
transform 1 0 304 0 -1 890
box -8 -3 16 105
use FILL  FILL_21
timestamp 1488311641
transform 1 0 312 0 -1 890
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_3
timestamp 1488311641
transform 1 0 362 0 1 790
box -7 -2 7 2
use $$M2_M1  $$M2_M1_8
timestamp 1488311641
transform 1 0 92 0 1 720
box -2 -2 2 2
use $$M2_M1  $$M2_M1_9
timestamp 1488311641
transform 1 0 132 0 1 731
box -2 -2 2 2
use $$M2_M1  $$M2_M1_10
timestamp 1488311641
transform 1 0 148 0 1 700
box -2 -2 2 2
use $$M3_M2  $$M3_M2_8
timestamp 1488311641
transform 1 0 148 0 1 700
box -3 -3 3 3
use $$M2_M1  $$M2_M1_11
timestamp 1488311641
transform 1 0 156 0 1 743
box -2 -2 2 2
use $$M3_M2  $$M3_M2_9
timestamp 1488311641
transform 1 0 180 0 1 720
box -3 -3 3 3
use $$M2_M1  $$M2_M1_12
timestamp 1488311641
transform 1 0 228 0 1 744
box -2 -2 2 2
use $$M2_M1  $$M2_M1_13
timestamp 1488311641
transform 1 0 212 0 1 731
box -2 -2 2 2
use $$M2_M1  $$M2_M1_14
timestamp 1488311641
transform 1 0 220 0 1 730
box -2 -2 2 2
use $$M3_M2  $$M3_M2_10
timestamp 1488311641
transform 1 0 220 0 1 730
box -3 -3 3 3
use $$M2_M1  $$M2_M1_15
timestamp 1488311641
transform 1 0 204 0 1 723
box -2 -2 2 2
use $$M3_M2  $$M3_M2_11
timestamp 1488311641
transform 1 0 228 0 1 720
box -3 -3 3 3
use $$M3_M2  $$M3_M2_12
timestamp 1488311641
transform 1 0 220 0 1 700
box -3 -3 3 3
use $$M2_M1  $$M2_M1_16
timestamp 1488311641
transform 1 0 252 0 1 724
box -2 -2 2 2
use $$M3_M2  $$M3_M2_13
timestamp 1488311641
transform 1 0 252 0 1 700
box -3 -3 3 3
use $$M3_M2  $$M3_M2_14
timestamp 1488311641
transform 1 0 316 0 1 730
box -3 -3 3 3
use $$M2_M1  $$M2_M1_17
timestamp 1488311641
transform 1 0 300 0 1 724
box -2 -2 2 2
use $$M2_M1  $$M2_M1_18
timestamp 1488311641
transform 1 0 316 0 1 721
box -2 -2 2 2
use $$M2_M1  $$M2_M1_19
timestamp 1488311641
transform 1 0 276 0 1 700
box -2 -2 2 2
use $$M2_M1  $$M2_M1_20
timestamp 1488311641
transform 1 0 308 0 1 700
box -2 -2 2 2
use $$M3_M2  $$M3_M2_15
timestamp 1488311641
transform 1 0 316 0 1 700
box -3 -3 3 3
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_4
timestamp 1488311641
transform 1 0 62 0 1 690
box -7 -2 7 2
use FILL  FILL_22
timestamp 1488311641
transform -1 0 88 0 1 690
box -8 -3 16 105
use FILL  FILL_23
timestamp 1488311641
transform -1 0 96 0 1 690
box -8 -3 16 105
use FILL  FILL_24
timestamp 1488311641
transform -1 0 104 0 1 690
box -8 -3 16 105
use $$M3_M2  $$M3_M2_16
timestamp 1488311641
transform 1 0 116 0 1 690
box -3 -3 3 3
use FILL  FILL_25
timestamp 1488311641
transform -1 0 112 0 1 690
box -8 -3 16 105
use FILL  FILL_26
timestamp 1488311641
transform -1 0 120 0 1 690
box -8 -3 16 105
use OAI21X1  OAI21X1_0
timestamp 1488311641
transform 1 0 120 0 1 690
box -8 -3 34 105
use FILL  FILL_27
timestamp 1488311641
transform -1 0 160 0 1 690
box -8 -3 16 105
use FILL  FILL_28
timestamp 1488311641
transform -1 0 168 0 1 690
box -8 -3 16 105
use FILL  FILL_29
timestamp 1488311641
transform -1 0 176 0 1 690
box -8 -3 16 105
use FILL  FILL_30
timestamp 1488311641
transform -1 0 184 0 1 690
box -8 -3 16 105
use FILL  FILL_31
timestamp 1488311641
transform -1 0 192 0 1 690
box -8 -3 16 105
use FILL  FILL_32
timestamp 1488311641
transform -1 0 200 0 1 690
box -8 -3 16 105
use $$M3_M2  $$M3_M2_17
timestamp 1488311641
transform 1 0 212 0 1 690
box -3 -3 3 3
use OAI21X1  OAI21X1_1
timestamp 1488311641
transform 1 0 200 0 1 690
box -8 -3 34 105
use FILL  FILL_33
timestamp 1488311641
transform -1 0 240 0 1 690
box -8 -3 16 105
use FILL  FILL_34
timestamp 1488311641
transform -1 0 248 0 1 690
box -8 -3 16 105
use $$M3_M2  $$M3_M2_18
timestamp 1488311641
transform 1 0 308 0 1 690
box -3 -3 3 3
use XOR2X1  XOR2X1_0
timestamp 1488311641
transform 1 0 248 0 1 690
box -8 -3 64 105
use INVX2  INVX2_2
timestamp 1488311641
transform -1 0 320 0 1 690
box -9 -3 26 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_5
timestamp 1488311641
transform 1 0 337 0 1 690
box -7 -2 7 2
use $$M2_M1  $$M2_M1_21
timestamp 1488311641
transform 1 0 108 0 1 680
box -2 -2 2 2
use $$M2_M1  $$M2_M1_22
timestamp 1488311641
transform 1 0 132 0 1 650
box -2 -2 2 2
use $$M2_M1  $$M2_M1_23
timestamp 1488311641
transform 1 0 124 0 1 643
box -2 -2 2 2
use $$M3_M2  $$M3_M2_19
timestamp 1488311641
transform 1 0 124 0 1 640
box -3 -3 3 3
use $$M2_M1  $$M2_M1_24
timestamp 1488311641
transform 1 0 108 0 1 630
box -2 -2 2 2
use $$M3_M2  $$M3_M2_20
timestamp 1488311641
transform 1 0 108 0 1 630
box -3 -3 3 3
use $$M3_M2  $$M3_M2_21
timestamp 1488311641
transform 1 0 204 0 1 670
box -3 -3 3 3
use $$M3_M2  $$M3_M2_22
timestamp 1488311641
transform 1 0 212 0 1 660
box -3 -3 3 3
use $$M2_M1  $$M2_M1_25
timestamp 1488311641
transform 1 0 188 0 1 650
box -2 -2 2 2
use $$M3_M2  $$M3_M2_23
timestamp 1488311641
transform 1 0 188 0 1 650
box -3 -3 3 3
use $$M2_M1  $$M2_M1_26
timestamp 1488311641
transform 1 0 204 0 1 653
box -2 -2 2 2
use $$M2_M1  $$M2_M1_27
timestamp 1488311641
transform 1 0 204 0 1 630
box -2 -2 2 2
use $$M2_M1  $$M2_M1_28
timestamp 1488311641
transform 1 0 228 0 1 650
box -2 -2 2 2
use $$M3_M2  $$M3_M2_24
timestamp 1488311641
transform 1 0 228 0 1 650
box -3 -3 3 3
use $$M2_M1  $$M2_M1_29
timestamp 1488311641
transform 1 0 228 0 1 640
box -2 -2 2 2
use $$M3_M2  $$M3_M2_25
timestamp 1488311641
transform 1 0 228 0 1 640
box -3 -3 3 3
use $$M2_M1  $$M2_M1_30
timestamp 1488311641
transform 1 0 236 0 1 630
box -2 -2 2 2
use $$M3_M2  $$M3_M2_26
timestamp 1488311641
transform 1 0 236 0 1 630
box -3 -3 3 3
use $$M3_M2  $$M3_M2_27
timestamp 1488311641
transform 1 0 284 0 1 660
box -3 -3 3 3
use $$M2_M1  $$M2_M1_31
timestamp 1488311641
transform 1 0 268 0 1 650
box -2 -2 2 2
use $$M2_M1  $$M2_M1_32
timestamp 1488311641
transform 1 0 284 0 1 649
box -2 -2 2 2
use $$M2_M1  $$M2_M1_33
timestamp 1488311641
transform 1 0 316 0 1 653
box -2 -2 2 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_6
timestamp 1488311641
transform 1 0 37 0 1 590
box -7 -2 7 2
use FILL  FILL_35
timestamp 1488311641
transform 1 0 80 0 -1 690
box -8 -3 16 105
use FILL  FILL_36
timestamp 1488311641
transform 1 0 88 0 -1 690
box -8 -3 16 105
use FILL  FILL_37
timestamp 1488311641
transform 1 0 96 0 -1 690
box -8 -3 16 105
use OAI21X1  OAI21X1_2
timestamp 1488311641
transform -1 0 136 0 -1 690
box -8 -3 34 105
use FILL  FILL_38
timestamp 1488311641
transform 1 0 136 0 -1 690
box -8 -3 16 105
use FILL  FILL_39
timestamp 1488311641
transform 1 0 144 0 -1 690
box -8 -3 16 105
use FILL  FILL_40
timestamp 1488311641
transform 1 0 152 0 -1 690
box -8 -3 16 105
use FILL  FILL_41
timestamp 1488311641
transform 1 0 160 0 -1 690
box -8 -3 16 105
use FILL  FILL_42
timestamp 1488311641
transform 1 0 168 0 -1 690
box -8 -3 16 105
use FILL  FILL_43
timestamp 1488311641
transform 1 0 176 0 -1 690
box -8 -3 16 105
use $$M3_M2  $$M3_M2_28
timestamp 1488311641
transform 1 0 204 0 1 590
box -3 -3 3 3
use INVX2  INVX2_3
timestamp 1488311641
transform -1 0 200 0 -1 690
box -9 -3 26 105
use $$M3_M2  $$M3_M2_29
timestamp 1488311641
transform 1 0 228 0 1 590
box -3 -3 3 3
use NAND2X1  NAND2X1_0
timestamp 1488311641
transform -1 0 224 0 -1 690
box -8 -3 32 105
use FILL  FILL_44
timestamp 1488311641
transform 1 0 224 0 -1 690
box -8 -3 16 105
use FILL  FILL_45
timestamp 1488311641
transform 1 0 232 0 -1 690
box -8 -3 16 105
use FILL  FILL_46
timestamp 1488311641
transform 1 0 240 0 -1 690
box -8 -3 16 105
use FILL  FILL_47
timestamp 1488311641
transform 1 0 248 0 -1 690
box -8 -3 16 105
use FILL  FILL_48
timestamp 1488311641
transform 1 0 256 0 -1 690
box -8 -3 16 105
use $$M3_M2  $$M3_M2_30
timestamp 1488311641
transform 1 0 300 0 1 590
box -3 -3 3 3
use OAI21X1  OAI21X1_3
timestamp 1488311641
transform -1 0 296 0 -1 690
box -8 -3 34 105
use FILL  FILL_49
timestamp 1488311641
transform 1 0 296 0 -1 690
box -8 -3 16 105
use FILL  FILL_50
timestamp 1488311641
transform 1 0 304 0 -1 690
box -8 -3 16 105
use FILL  FILL_51
timestamp 1488311641
transform 1 0 312 0 -1 690
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_7
timestamp 1488311641
transform 1 0 362 0 1 590
box -7 -2 7 2
use $$M3_M2  $$M3_M2_31
timestamp 1488311641
transform 1 0 92 0 1 500
box -3 -3 3 3
use $$M2_M1  $$M2_M1_34
timestamp 1488311641
transform 1 0 108 0 1 580
box -2 -2 2 2
use $$M3_M2  $$M3_M2_32
timestamp 1488311641
transform 1 0 108 0 1 580
box -3 -3 3 3
use $$M3_M2  $$M3_M2_33
timestamp 1488311641
transform 1 0 132 0 1 580
box -3 -3 3 3
use $$M2_M1  $$M2_M1_35
timestamp 1488311641
transform 1 0 132 0 1 520
box -2 -2 2 2
use $$M3_M2  $$M3_M2_34
timestamp 1488311641
transform 1 0 132 0 1 520
box -3 -3 3 3
use $$M2_M1  $$M2_M1_36
timestamp 1488311641
transform 1 0 140 0 1 511
box -2 -2 2 2
use $$M3_M2  $$M3_M2_35
timestamp 1488311641
transform 1 0 124 0 1 500
box -3 -3 3 3
use $$M3_M2  $$M3_M2_36
timestamp 1488311641
transform 1 0 172 0 1 530
box -3 -3 3 3
use $$M2_M1  $$M2_M1_37
timestamp 1488311641
transform 1 0 188 0 1 550
box -2 -2 2 2
use $$M2_M1  $$M2_M1_38
timestamp 1488311641
transform 1 0 196 0 1 500
box -2 -2 2 2
use $$M2_M1  $$M2_M1_39
timestamp 1488311641
transform 1 0 220 0 1 520
box -2 -2 2 2
use $$M3_M2  $$M3_M2_37
timestamp 1488311641
transform 1 0 220 0 1 520
box -3 -3 3 3
use $$M2_M1  $$M2_M1_40
timestamp 1488311641
transform 1 0 236 0 1 530
box -2 -2 2 2
use $$M3_M2  $$M3_M2_38
timestamp 1488311641
transform 1 0 236 0 1 530
box -3 -3 3 3
use $$M2_M1  $$M2_M1_41
timestamp 1488311641
transform 1 0 292 0 1 530
box -2 -2 2 2
use $$M2_M1  $$M2_M1_42
timestamp 1488311641
transform 1 0 300 0 1 530
box -2 -2 2 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_8
timestamp 1488311641
transform 1 0 62 0 1 490
box -7 -2 7 2
use FILL  FILL_52
timestamp 1488311641
transform -1 0 88 0 1 490
box -8 -3 16 105
use FILL  FILL_53
timestamp 1488311641
transform -1 0 96 0 1 490
box -8 -3 16 105
use FILL  FILL_54
timestamp 1488311641
transform -1 0 104 0 1 490
box -8 -3 16 105
use FILL  FILL_55
timestamp 1488311641
transform -1 0 112 0 1 490
box -8 -3 16 105
use OR2X1  OR2X1_0
timestamp 1488311641
transform -1 0 144 0 1 490
box -8 -3 40 105
use FILL  FILL_56
timestamp 1488311641
transform -1 0 152 0 1 490
box -8 -3 16 105
use FILL  FILL_57
timestamp 1488311641
transform -1 0 160 0 1 490
box -8 -3 16 105
use FILL  FILL_58
timestamp 1488311641
transform -1 0 168 0 1 490
box -8 -3 16 105
use FILL  FILL_59
timestamp 1488311641
transform -1 0 176 0 1 490
box -8 -3 16 105
use FILL  FILL_60
timestamp 1488311641
transform -1 0 184 0 1 490
box -8 -3 16 105
use FILL  FILL_61
timestamp 1488311641
transform -1 0 192 0 1 490
box -8 -3 16 105
use NAND2X1  NAND2X1_1
timestamp 1488311641
transform -1 0 216 0 1 490
box -8 -3 32 105
use FILL  FILL_62
timestamp 1488311641
transform -1 0 224 0 1 490
box -8 -3 16 105
use FILL  FILL_63
timestamp 1488311641
transform -1 0 232 0 1 490
box -8 -3 16 105
use FILL  FILL_64
timestamp 1488311641
transform -1 0 240 0 1 490
box -8 -3 16 105
use FILL  FILL_65
timestamp 1488311641
transform -1 0 248 0 1 490
box -8 -3 16 105
use FILL  FILL_66
timestamp 1488311641
transform -1 0 256 0 1 490
box -8 -3 16 105
use $$M3_M2  $$M3_M2_39
timestamp 1488311641
transform 1 0 268 0 1 490
box -3 -3 3 3
use FILL  FILL_67
timestamp 1488311641
transform -1 0 264 0 1 490
box -8 -3 16 105
use FILL  FILL_68
timestamp 1488311641
transform -1 0 272 0 1 490
box -8 -3 16 105
use $$M3_M2  $$M3_M2_40
timestamp 1488311641
transform 1 0 300 0 1 490
box -3 -3 3 3
use AND2X2  AND2X2_0
timestamp 1488311641
transform -1 0 304 0 1 490
box -8 -3 40 105
use FILL  FILL_69
timestamp 1488311641
transform -1 0 312 0 1 490
box -8 -3 16 105
use FILL  FILL_70
timestamp 1488311641
transform -1 0 320 0 1 490
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_9
timestamp 1488311641
transform 1 0 337 0 1 490
box -7 -2 7 2
use $$M2_M1  $$M2_M1_43
timestamp 1488311641
transform 1 0 92 0 1 480
box -2 -2 2 2
use $$M3_M2  $$M3_M2_41
timestamp 1488311641
transform 1 0 92 0 1 480
box -3 -3 3 3
use $$M2_M1  $$M2_M1_44
timestamp 1488311641
transform 1 0 124 0 1 453
box -2 -2 2 2
use $$M3_M2  $$M3_M2_42
timestamp 1488311641
transform 1 0 140 0 1 470
box -3 -3 3 3
use $$M3_M2  $$M3_M2_43
timestamp 1488311641
transform 1 0 164 0 1 480
box -3 -3 3 3
use $$M2_M1  $$M2_M1_45
timestamp 1488311641
transform 1 0 164 0 1 450
box -2 -2 2 2
use $$M2_M1  $$M2_M1_46
timestamp 1488311641
transform 1 0 204 0 1 440
box -2 -2 2 2
use $$M3_M2  $$M3_M2_44
timestamp 1488311641
transform 1 0 204 0 1 440
box -3 -3 3 3
use $$M2_M1  $$M2_M1_47
timestamp 1488311641
transform 1 0 220 0 1 430
box -2 -2 2 2
use $$M2_M1  $$M2_M1_48
timestamp 1488311641
transform 1 0 252 0 1 453
box -2 -2 2 2
use $$M3_M2  $$M3_M2_45
timestamp 1488311641
transform 1 0 244 0 1 440
box -3 -3 3 3
use $$M3_M2  $$M3_M2_46
timestamp 1488311641
transform 1 0 260 0 1 430
box -3 -3 3 3
use $$M2_M1  $$M2_M1_49
timestamp 1488311641
transform 1 0 260 0 1 400
box -2 -2 2 2
use $$M2_M1  $$M2_M1_50
timestamp 1488311641
transform 1 0 284 0 1 449
box -2 -2 2 2
use $$M2_M1  $$M2_M1_51
timestamp 1488311641
transform 1 0 289 0 1 400
box -2 -2 2 2
use $$M2_M1  $$M2_M1_52
timestamp 1488311641
transform 1 0 308 0 1 430
box -2 -2 2 2
use $$M3_M2  $$M3_M2_47
timestamp 1488311641
transform 1 0 308 0 1 430
box -3 -3 3 3
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_10
timestamp 1488311641
transform 1 0 37 0 1 390
box -7 -2 7 2
use FILL  FILL_71
timestamp 1488311641
transform 1 0 80 0 -1 490
box -8 -3 16 105
use FILL  FILL_72
timestamp 1488311641
transform 1 0 88 0 -1 490
box -8 -3 16 105
use INVX2  INVX2_4
timestamp 1488311641
transform -1 0 112 0 -1 490
box -9 -3 26 105
use FILL  FILL_73
timestamp 1488311641
transform 1 0 112 0 -1 490
box -8 -3 16 105
use FILL  FILL_74
timestamp 1488311641
transform 1 0 120 0 -1 490
box -8 -3 16 105
use FILL  FILL_75
timestamp 1488311641
transform 1 0 128 0 -1 490
box -8 -3 16 105
use FILL  FILL_76
timestamp 1488311641
transform 1 0 136 0 -1 490
box -8 -3 16 105
use FILL  FILL_77
timestamp 1488311641
transform 1 0 144 0 -1 490
box -8 -3 16 105
use FILL  FILL_78
timestamp 1488311641
transform 1 0 152 0 -1 490
box -8 -3 16 105
use FILL  FILL_79
timestamp 1488311641
transform 1 0 160 0 -1 490
box -8 -3 16 105
use FILL  FILL_80
timestamp 1488311641
transform 1 0 168 0 -1 490
box -8 -3 16 105
use FILL  FILL_81
timestamp 1488311641
transform 1 0 176 0 -1 490
box -8 -3 16 105
use FILL  FILL_82
timestamp 1488311641
transform 1 0 184 0 -1 490
box -8 -3 16 105
use FILL  FILL_83
timestamp 1488311641
transform 1 0 192 0 -1 490
box -8 -3 16 105
use FILL  FILL_84
timestamp 1488311641
transform 1 0 200 0 -1 490
box -8 -3 16 105
use NAND3X1  NAND3X1_0
timestamp 1488311641
transform 1 0 208 0 -1 490
box -8 -3 40 105
use FILL  FILL_85
timestamp 1488311641
transform 1 0 240 0 -1 490
box -8 -3 16 105
use FILL  FILL_86
timestamp 1488311641
transform 1 0 248 0 -1 490
box -8 -3 16 105
use FILL  FILL_87
timestamp 1488311641
transform 1 0 256 0 -1 490
box -8 -3 16 105
use FILL  FILL_88
timestamp 1488311641
transform 1 0 264 0 -1 490
box -8 -3 16 105
use OAI21X1  OAI21X1_4
timestamp 1488311641
transform 1 0 272 0 -1 490
box -8 -3 34 105
use FILL  FILL_89
timestamp 1488311641
transform 1 0 304 0 -1 490
box -8 -3 16 105
use FILL  FILL_90
timestamp 1488311641
transform 1 0 312 0 -1 490
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_11
timestamp 1488311641
transform 1 0 362 0 1 390
box -7 -2 7 2
use $$M2_M1  $$M2_M1_53
timestamp 1488311641
transform 1 0 108 0 1 340
box -2 -2 2 2
use $$M3_M2  $$M3_M2_48
timestamp 1488311641
transform 1 0 108 0 1 340
box -3 -3 3 3
use $$M2_M1  $$M2_M1_54
timestamp 1488311641
transform 1 0 92 0 1 321
box -2 -2 2 2
use $$M3_M2  $$M3_M2_49
timestamp 1488311641
transform 1 0 92 0 1 320
box -3 -3 3 3
use $$M2_M1  $$M2_M1_55
timestamp 1488311641
transform 1 0 108 0 1 323
box -2 -2 2 2
use $$M3_M2  $$M3_M2_50
timestamp 1488311641
transform 1 0 108 0 1 320
box -3 -3 3 3
use $$M3_M2  $$M3_M2_51
timestamp 1488311641
transform 1 0 124 0 1 370
box -3 -3 3 3
use $$M2_M1  $$M2_M1_56
timestamp 1488311641
transform 1 0 124 0 1 350
box -2 -2 2 2
use $$M3_M2  $$M3_M2_52
timestamp 1488311641
transform 1 0 124 0 1 340
box -3 -3 3 3
use $$M2_M1  $$M2_M1_57
timestamp 1488311641
transform 1 0 132 0 1 300
box -2 -2 2 2
use $$M2_M1  $$M2_M1_58
timestamp 1488311641
transform 1 0 180 0 1 380
box -2 -2 2 2
use $$M3_M2  $$M3_M2_53
timestamp 1488311641
transform 1 0 180 0 1 370
box -3 -3 3 3
use $$M2_M1  $$M2_M1_59
timestamp 1488311641
transform 1 0 172 0 1 350
box -2 -2 2 2
use $$M2_M1  $$M2_M1_60
timestamp 1488311641
transform 1 0 188 0 1 340
box -2 -2 2 2
use $$M3_M2  $$M3_M2_54
timestamp 1488311641
transform 1 0 172 0 1 330
box -3 -3 3 3
use $$M2_M1  $$M2_M1_61
timestamp 1488311641
transform 1 0 180 0 1 333
box -2 -2 2 2
use $$M3_M2  $$M3_M2_55
timestamp 1488311641
transform 1 0 220 0 1 330
box -3 -3 3 3
use $$M2_M1  $$M2_M1_62
timestamp 1488311641
transform 1 0 220 0 1 323
box -2 -2 2 2
use $$M3_M2  $$M3_M2_56
timestamp 1488311641
transform 1 0 228 0 1 320
box -3 -3 3 3
use $$M2_M1  $$M2_M1_63
timestamp 1488311641
transform 1 0 260 0 1 350
box -2 -2 2 2
use $$M3_M2  $$M3_M2_57
timestamp 1488311641
transform 1 0 244 0 1 340
box -3 -3 3 3
use $$M2_M1  $$M2_M1_64
timestamp 1488311641
transform 1 0 244 0 1 337
box -2 -2 2 2
use $$M2_M1  $$M2_M1_65
timestamp 1488311641
transform 1 0 260 0 1 320
box -2 -2 2 2
use $$M3_M2  $$M3_M2_58
timestamp 1488311641
transform 1 0 260 0 1 320
box -3 -3 3 3
use $$M2_M1  $$M2_M1_66
timestamp 1488311641
transform 1 0 316 0 1 380
box -2 -2 2 2
use $$M2_M1  $$M2_M1_67
timestamp 1488311641
transform 1 0 308 0 1 321
box -2 -2 2 2
use $$M3_M2  $$M3_M2_59
timestamp 1488311641
transform 1 0 308 0 1 320
box -3 -3 3 3
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_12
timestamp 1488311641
transform 1 0 62 0 1 290
box -7 -2 7 2
use FILL  FILL_91
timestamp 1488311641
transform -1 0 88 0 1 290
box -8 -3 16 105
use INVX2  INVX2_5
timestamp 1488311641
transform 1 0 88 0 1 290
box -9 -3 26 105
use NAND2X1  NAND2X1_2
timestamp 1488311641
transform 1 0 104 0 1 290
box -8 -3 32 105
use FILL  FILL_92
timestamp 1488311641
transform -1 0 136 0 1 290
box -8 -3 16 105
use FILL  FILL_93
timestamp 1488311641
transform -1 0 144 0 1 290
box -8 -3 16 105
use FILL  FILL_94
timestamp 1488311641
transform -1 0 152 0 1 290
box -8 -3 16 105
use FILL  FILL_95
timestamp 1488311641
transform -1 0 160 0 1 290
box -8 -3 16 105
use NAND3X1  NAND3X1_1
timestamp 1488311641
transform -1 0 192 0 1 290
box -8 -3 40 105
use FILL  FILL_96
timestamp 1488311641
transform -1 0 200 0 1 290
box -8 -3 16 105
use $$M3_M2  $$M3_M2_60
timestamp 1488311641
transform 1 0 212 0 1 290
box -3 -3 3 3
use FILL  FILL_97
timestamp 1488311641
transform -1 0 208 0 1 290
box -8 -3 16 105
use FILL  FILL_98
timestamp 1488311641
transform -1 0 216 0 1 290
box -8 -3 16 105
use FILL  FILL_99
timestamp 1488311641
transform -1 0 224 0 1 290
box -8 -3 16 105
use FILL  FILL_100
timestamp 1488311641
transform -1 0 232 0 1 290
box -8 -3 16 105
use OAI21X1  OAI21X1_5
timestamp 1488311641
transform 1 0 232 0 1 290
box -8 -3 34 105
use FILL  FILL_101
timestamp 1488311641
transform -1 0 272 0 1 290
box -8 -3 16 105
use FILL  FILL_102
timestamp 1488311641
transform -1 0 280 0 1 290
box -8 -3 16 105
use FILL  FILL_103
timestamp 1488311641
transform -1 0 288 0 1 290
box -8 -3 16 105
use FILL  FILL_104
timestamp 1488311641
transform -1 0 296 0 1 290
box -8 -3 16 105
use FILL  FILL_105
timestamp 1488311641
transform -1 0 304 0 1 290
box -8 -3 16 105
use INVX2  INVX2_6
timestamp 1488311641
transform 1 0 304 0 1 290
box -9 -3 26 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_13
timestamp 1488311641
transform 1 0 337 0 1 290
box -7 -2 7 2
use $$M3_M2  $$M3_M2_61
timestamp 1488311641
transform 1 0 20 0 1 260
box -3 -3 3 3
use $$M3_M2  $$M3_M2_62
timestamp 1488311641
transform 1 0 100 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_68
timestamp 1488311641
transform 1 0 100 0 1 253
box -2 -2 2 2
use $$M3_M2  $$M3_M2_63
timestamp 1488311641
transform 1 0 124 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_69
timestamp 1488311641
transform 1 0 116 0 1 230
box -2 -2 2 2
use $$M2_M1  $$M2_M1_70
timestamp 1488311641
transform 1 0 108 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_64
timestamp 1488311641
transform 1 0 140 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_71
timestamp 1488311641
transform 1 0 156 0 1 280
box -2 -2 2 2
use $$M2_M1  $$M2_M1_72
timestamp 1488311641
transform 1 0 148 0 1 250
box -2 -2 2 2
use $$M3_M2  $$M3_M2_65
timestamp 1488311641
transform 1 0 180 0 1 280
box -3 -3 3 3
use $$M2_M1  $$M2_M1_73
timestamp 1488311641
transform 1 0 172 0 1 247
box -2 -2 2 2
use $$M2_M1  $$M2_M1_74
timestamp 1488311641
transform 1 0 180 0 1 240
box -2 -2 2 2
use $$M2_M1  $$M2_M1_75
timestamp 1488311641
transform 1 0 164 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_66
timestamp 1488311641
transform 1 0 164 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_76
timestamp 1488311641
transform 1 0 204 0 1 280
box -2 -2 2 2
use $$M3_M2  $$M3_M2_67
timestamp 1488311641
transform 1 0 204 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_77
timestamp 1488311641
transform 1 0 204 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_68
timestamp 1488311641
transform 1 0 228 0 1 280
box -3 -3 3 3
use $$M2_M1  $$M2_M1_78
timestamp 1488311641
transform 1 0 252 0 1 270
box -2 -2 2 2
use $$M3_M2  $$M3_M2_69
timestamp 1488311641
transform 1 0 252 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_70
timestamp 1488311641
transform 1 0 220 0 1 260
box -3 -3 3 3
use $$M3_M2  $$M3_M2_71
timestamp 1488311641
transform 1 0 244 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_79
timestamp 1488311641
transform 1 0 220 0 1 256
box -2 -2 2 2
use $$M2_M1  $$M2_M1_80
timestamp 1488311641
transform 1 0 228 0 1 253
box -2 -2 2 2
use $$M3_M2  $$M3_M2_72
timestamp 1488311641
transform 1 0 236 0 1 250
box -3 -3 3 3
use $$M3_M2  $$M3_M2_73
timestamp 1488311641
transform 1 0 228 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_81
timestamp 1488311641
transform 1 0 236 0 1 243
box -2 -2 2 2
use $$M3_M2  $$M3_M2_74
timestamp 1488311641
transform 1 0 244 0 1 230
box -3 -3 3 3
use $$M3_M2  $$M3_M2_75
timestamp 1488311641
transform 1 0 276 0 1 260
box -3 -3 3 3
use $$M2_M1  $$M2_M1_82
timestamp 1488311641
transform 1 0 276 0 1 255
box -2 -2 2 2
use $$M2_M1  $$M2_M1_83
timestamp 1488311641
transform 1 0 268 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_76
timestamp 1488311641
transform 1 0 268 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_84
timestamp 1488311641
transform 1 0 284 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_77
timestamp 1488311641
transform 1 0 284 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_85
timestamp 1488311641
transform 1 0 292 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_78
timestamp 1488311641
transform 1 0 308 0 1 260
box -3 -3 3 3
use $$M3_M2  $$M3_M2_79
timestamp 1488311641
transform 1 0 316 0 1 240
box -3 -3 3 3
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_14
timestamp 1488311641
transform 1 0 37 0 1 190
box -7 -2 7 2
use FILL  FILL_106
timestamp 1488311641
transform 1 0 80 0 -1 290
box -8 -3 16 105
use FILL  FILL_107
timestamp 1488311641
transform 1 0 88 0 -1 290
box -8 -3 16 105
use NAND2X1  NAND2X1_3
timestamp 1488311641
transform 1 0 96 0 -1 290
box -8 -3 32 105
use FILL  FILL_108
timestamp 1488311641
transform 1 0 120 0 -1 290
box -8 -3 16 105
use FILL  FILL_109
timestamp 1488311641
transform 1 0 128 0 -1 290
box -8 -3 16 105
use FILL  FILL_110
timestamp 1488311641
transform 1 0 136 0 -1 290
box -8 -3 16 105
use FILL  FILL_111
timestamp 1488311641
transform 1 0 144 0 -1 290
box -8 -3 16 105
use NAND3X1  NAND3X1_2
timestamp 1488311641
transform -1 0 184 0 -1 290
box -8 -3 40 105
use FILL  FILL_112
timestamp 1488311641
transform 1 0 184 0 -1 290
box -8 -3 16 105
use FILL  FILL_113
timestamp 1488311641
transform 1 0 192 0 -1 290
box -8 -3 16 105
use NAND2X1  NAND2X1_4
timestamp 1488311641
transform -1 0 224 0 -1 290
box -8 -3 32 105
use OAI21X1  OAI21X1_6
timestamp 1488311641
transform 1 0 224 0 -1 290
box -8 -3 34 105
use FILL  FILL_114
timestamp 1488311641
transform 1 0 256 0 -1 290
box -8 -3 16 105
use FILL  FILL_115
timestamp 1488311641
transform 1 0 264 0 -1 290
box -8 -3 16 105
use NAND2X1  NAND2X1_5
timestamp 1488311641
transform 1 0 272 0 -1 290
box -8 -3 32 105
use FILL  FILL_116
timestamp 1488311641
transform 1 0 296 0 -1 290
box -8 -3 16 105
use FILL  FILL_117
timestamp 1488311641
transform 1 0 304 0 -1 290
box -8 -3 16 105
use FILL  FILL_118
timestamp 1488311641
transform 1 0 312 0 -1 290
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_15
timestamp 1488311641
transform 1 0 362 0 1 190
box -7 -2 7 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_16
timestamp 1488311641
transform 1 0 62 0 1 90
box -7 -2 7 2
use FILL  FILL_119
timestamp 1488311641
transform -1 0 88 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_86
timestamp 1488311641
transform 1 0 100 0 1 147
box -2 -2 2 2
use FILL  FILL_120
timestamp 1488311641
transform -1 0 96 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_80
timestamp 1488311641
transform 1 0 108 0 1 160
box -3 -3 3 3
use $$M3_M2  $$M3_M2_81
timestamp 1488311641
transform 1 0 124 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_87
timestamp 1488311641
transform 1 0 124 0 1 137
box -2 -2 2 2
use $$M2_M1  $$M2_M1_88
timestamp 1488311641
transform 1 0 108 0 1 100
box -2 -2 2 2
use FILL  FILL_121
timestamp 1488311641
transform -1 0 104 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_89
timestamp 1488311641
transform 1 0 132 0 1 127
box -2 -2 2 2
use OAI21X1  OAI21X1_7
timestamp 1488311641
transform -1 0 136 0 1 90
box -8 -3 34 105
use FILL  FILL_122
timestamp 1488311641
transform -1 0 144 0 1 90
box -8 -3 16 105
use FILL  FILL_123
timestamp 1488311641
transform -1 0 152 0 1 90
box -8 -3 16 105
use FILL  FILL_124
timestamp 1488311641
transform -1 0 160 0 1 90
box -8 -3 16 105
use FILL  FILL_125
timestamp 1488311641
transform -1 0 168 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_90
timestamp 1488311641
transform 1 0 188 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_82
timestamp 1488311641
transform 1 0 180 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_91
timestamp 1488311641
transform 1 0 180 0 1 117
box -2 -2 2 2
use FILL  FILL_126
timestamp 1488311641
transform -1 0 176 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_83
timestamp 1488311641
transform 1 0 196 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_92
timestamp 1488311641
transform 1 0 196 0 1 133
box -2 -2 2 2
use $$M3_M2  $$M3_M2_84
timestamp 1488311641
transform 1 0 196 0 1 130
box -3 -3 3 3
use NOR2X1  NOR2X1_0
timestamp 1488311641
transform 1 0 176 0 1 90
box -8 -3 32 105
use $$M2_M1  $$M2_M1_93
timestamp 1488311641
transform 1 0 212 0 1 117
box -2 -2 2 2
use FILL  FILL_127
timestamp 1488311641
transform -1 0 208 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_94
timestamp 1488311641
transform 1 0 228 0 1 139
box -2 -2 2 2
use NOR2X1  NOR2X1_1
timestamp 1488311641
transform 1 0 208 0 1 90
box -8 -3 32 105
use FILL  FILL_128
timestamp 1488311641
transform -1 0 240 0 1 90
box -8 -3 16 105
use FILL  FILL_129
timestamp 1488311641
transform -1 0 248 0 1 90
box -8 -3 16 105
use FILL  FILL_130
timestamp 1488311641
transform -1 0 256 0 1 90
box -8 -3 16 105
use FILL  FILL_131
timestamp 1488311641
transform -1 0 264 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_95
timestamp 1488311641
transform 1 0 284 0 1 150
box -2 -2 2 2
use $$M2_M1  $$M2_M1_96
timestamp 1488311641
transform 1 0 276 0 1 130
box -2 -2 2 2
use $$M3_M2  $$M3_M2_85
timestamp 1488311641
transform 1 0 276 0 1 130
box -3 -3 3 3
use $$M3_M2  $$M3_M2_86
timestamp 1488311641
transform 1 0 276 0 1 120
box -3 -3 3 3
use $$M3_M2  $$M3_M2_87
timestamp 1488311641
transform 1 0 292 0 1 120
box -3 -3 3 3
use $$M2_M1  $$M2_M1_97
timestamp 1488311641
transform 1 0 292 0 1 117
box -2 -2 2 2
use NAND2X1  NAND2X1_6
timestamp 1488311641
transform 1 0 264 0 1 90
box -8 -3 32 105
use $$M2_M1  $$M2_M1_98
timestamp 1488311641
transform 1 0 308 0 1 180
box -2 -2 2 2
use $$M2_M1  $$M2_M1_99
timestamp 1488311641
transform 1 0 308 0 1 130
box -2 -2 2 2
use NOR2X1  NOR2X1_2
timestamp 1488311641
transform 1 0 288 0 1 90
box -8 -3 32 105
use FILL  FILL_132
timestamp 1488311641
transform -1 0 320 0 1 90
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_17
timestamp 1488311641
transform 1 0 337 0 1 90
box -7 -2 7 2
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_4
timestamp 1488311641
transform 1 0 62 0 1 72
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_5
timestamp 1488311641
transform 1 0 337 0 1 72
box -7 -7 7 7
use $$M3_M2  $$M3_M2_88
timestamp 1488311641
transform 1 0 108 0 1 60
box -3 -3 3 3
use $$M3_M2  $$M3_M2_89
timestamp 1488311641
transform 1 0 284 0 1 60
box -3 -3 3 3
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_6
timestamp 1488311641
transform 1 0 37 0 1 47
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_7
timestamp 1488311641
transform 1 0 362 0 1 47
box -7 -7 7 7
<< labels >>
flabel metal3 2 470 2 470 4 FreeSans 26 0 0 0 alu_op[0]
flabel metal3 2 920 2 920 4 FreeSans 26 0 0 0 op[2]
flabel metal3 2 700 2 700 4 FreeSans 26 0 0 0 op[3]
flabel metal3 2 490 2 490 4 FreeSans 26 0 0 0 op[4]
flabel metal3 2 270 2 270 4 FreeSans 26 0 0 0 op[5]
flabel metal3 2 60 2 60 4 FreeSans 26 0 0 0 op[6]
flabel metal2 44 978 44 978 4 FreeSans 26 0 0 0 op[1]
flabel metal2 356 978 356 978 4 FreeSans 26 0 0 0 op[0]
flabel metal3 397 700 397 700 4 FreeSans 26 0 0 0 funct[2]
flabel metal3 397 490 397 490 4 FreeSans 26 0 0 0 funct[3]
flabel metal3 397 920 397 920 4 FreeSans 26 0 0 0 funct[1]
flabel metal3 397 270 397 270 4 FreeSans 26 0 0 0 funct[4]
flabel metal3 397 60 397 60 4 FreeSans 26 0 0 0 funct[5]
flabel metal2 44 1 44 1 4 FreeSans 26 0 0 0 funct[0]
flabel metal2 356 1 356 1 4 FreeSans 26 0 0 0 alu_op[1]
<< end >>
                                                                                                                                                                                                                                                                             alu.mag                                                                                             0000644 �    Asz0000145 00000060655 13045425605 010263  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1486236549
<< nwell >>
rect 124 175 125 178
<< metal1 >>
rect 30 856 294 864
rect 348 803 352 807
rect -2 746 294 754
rect -2 662 366 664
rect -2 658 360 662
rect 364 658 366 662
rect -2 656 366 658
rect -2 636 294 644
rect -2 552 366 554
rect -2 548 360 552
rect 364 548 366 552
rect -2 546 366 548
rect -2 526 294 534
rect -2 442 366 444
rect -2 438 360 442
rect 364 438 366 442
rect -2 436 366 438
rect -2 416 294 424
rect -2 332 366 334
rect -2 328 360 332
rect 364 328 366 332
rect -2 326 366 328
rect -2 306 294 314
rect -2 222 366 224
rect -2 218 360 222
rect 364 218 366 222
rect -2 216 366 218
rect -2 196 294 204
rect -2 112 366 114
rect -2 108 360 112
rect 364 108 366 112
rect -2 106 366 108
rect -2 86 294 94
rect 356 33 363 37
rect -2 -4 294 4
<< m2contact >>
rect 344 803 348 807
rect 352 803 356 807
rect 360 768 364 772
rect 360 658 364 662
rect 360 548 364 552
rect 360 438 364 442
rect 360 328 364 332
rect 360 218 364 222
rect 360 108 364 112
rect 352 33 356 37
<< metal2 >>
rect 47 922 53 923
rect 47 918 48 922
rect 52 918 53 922
rect 47 917 53 918
rect 191 922 197 923
rect 191 918 192 922
rect 196 918 197 922
rect 288 918 292 922
rect 320 918 324 922
rect 191 917 197 918
rect 111 852 117 853
rect 111 848 112 852
rect 116 848 117 852
rect 111 847 117 848
rect 143 852 149 853
rect 143 848 144 852
rect 148 848 149 852
rect 143 847 149 848
rect 159 852 165 853
rect 159 848 160 852
rect 164 848 165 852
rect 159 847 165 848
rect 31 842 37 843
rect 31 838 32 842
rect 36 838 37 842
rect 31 837 37 838
rect 95 822 101 823
rect 95 818 96 822
rect 100 818 101 822
rect 95 817 101 818
rect 87 812 93 813
rect 87 808 88 812
rect 92 808 93 812
rect 96 809 100 817
rect 87 807 93 808
rect 112 801 116 847
rect 119 842 125 843
rect 119 838 120 842
rect 124 838 125 842
rect 119 837 125 838
rect 120 832 125 837
rect 144 818 148 847
rect 151 842 157 843
rect 151 838 152 842
rect 156 838 157 842
rect 151 837 157 838
rect 128 803 132 811
rect 127 802 133 803
rect 127 798 128 802
rect 132 798 133 802
rect 127 797 133 798
rect 152 793 156 837
rect 160 803 164 847
rect 167 812 173 813
rect 167 808 168 812
rect 172 808 173 812
rect 167 807 173 808
rect 15 782 21 783
rect 15 778 16 782
rect 20 778 21 782
rect 15 777 21 778
rect 0 673 4 706
rect 16 687 20 777
rect 111 742 117 743
rect 111 738 112 742
rect 116 738 117 742
rect 111 737 117 738
rect 143 742 149 743
rect 143 738 144 742
rect 148 738 149 742
rect 143 737 149 738
rect 159 742 165 743
rect 159 738 160 742
rect 164 738 165 742
rect 159 737 165 738
rect 31 732 37 733
rect 31 728 32 732
rect 36 728 37 732
rect 31 727 37 728
rect 95 712 101 713
rect 95 708 96 712
rect 100 708 101 712
rect 95 707 101 708
rect 87 702 93 703
rect 87 698 88 702
rect 92 698 93 702
rect 96 699 100 707
rect 87 697 93 698
rect 112 691 116 737
rect 119 732 125 733
rect 119 728 120 732
rect 124 728 125 732
rect 119 727 125 728
rect 120 722 125 727
rect 144 708 148 737
rect 151 732 157 733
rect 151 728 152 732
rect 156 728 157 732
rect 151 727 157 728
rect 128 693 132 701
rect 127 692 133 693
rect 127 688 128 692
rect 132 688 133 692
rect 127 687 133 688
rect 152 683 156 727
rect 160 693 164 737
rect 167 702 173 703
rect 167 698 168 702
rect 172 698 173 702
rect 167 697 173 698
rect -1 672 5 673
rect -1 668 0 672
rect 4 668 5 672
rect -1 667 5 668
rect 111 632 117 633
rect 111 628 112 632
rect 116 628 117 632
rect 111 627 117 628
rect 143 632 149 633
rect 143 628 144 632
rect 148 628 149 632
rect 143 627 149 628
rect 159 632 165 633
rect 159 628 160 632
rect 164 628 165 632
rect 159 627 165 628
rect 31 622 37 623
rect 31 618 32 622
rect 36 618 37 622
rect 31 617 37 618
rect 95 602 101 603
rect 95 598 96 602
rect 100 598 101 602
rect 95 597 101 598
rect 87 592 93 593
rect 87 588 88 592
rect 92 588 93 592
rect 96 589 100 597
rect 87 587 93 588
rect 112 581 116 627
rect 119 622 125 623
rect 119 618 120 622
rect 124 618 125 622
rect 119 617 125 618
rect 120 612 125 617
rect 144 598 148 627
rect 151 622 157 623
rect 151 618 152 622
rect 156 618 157 622
rect 151 617 157 618
rect 128 583 132 591
rect 127 582 133 583
rect 127 578 128 582
rect 132 578 133 582
rect 127 577 133 578
rect 152 573 156 617
rect 160 583 164 627
rect 167 592 173 593
rect 167 588 168 592
rect 172 588 173 592
rect 167 587 173 588
rect -1 562 5 563
rect -1 558 0 562
rect 4 558 5 562
rect -1 557 5 558
rect 0 484 4 557
rect 111 522 117 523
rect 111 518 112 522
rect 116 518 117 522
rect 111 517 117 518
rect 143 522 149 523
rect 143 518 144 522
rect 148 518 149 522
rect 143 517 149 518
rect 159 522 165 523
rect 159 518 160 522
rect 164 518 165 522
rect 159 517 165 518
rect 31 512 37 513
rect 31 508 32 512
rect 36 508 37 512
rect 31 507 37 508
rect 95 492 101 493
rect 95 488 96 492
rect 100 488 101 492
rect 95 487 101 488
rect 87 482 93 483
rect 87 478 88 482
rect 92 478 93 482
rect 96 479 100 487
rect 87 477 93 478
rect 112 471 116 517
rect 119 512 125 513
rect 119 508 120 512
rect 124 508 125 512
rect 119 507 125 508
rect 120 502 125 507
rect 144 488 148 517
rect 151 512 157 513
rect 151 508 152 512
rect 156 508 157 512
rect 151 507 157 508
rect 128 473 132 481
rect 127 472 133 473
rect 16 453 20 469
rect 127 468 128 472
rect 132 468 133 472
rect 127 467 133 468
rect 152 463 156 507
rect 160 473 164 517
rect 167 482 173 483
rect 167 478 168 482
rect 172 478 173 482
rect 167 477 173 478
rect 15 452 21 453
rect 15 448 16 452
rect 20 448 21 452
rect 15 447 21 448
rect 111 412 117 413
rect 111 408 112 412
rect 116 408 117 412
rect 111 407 117 408
rect 143 412 149 413
rect 143 408 144 412
rect 148 408 149 412
rect 143 407 149 408
rect 159 412 165 413
rect 159 408 160 412
rect 164 408 165 412
rect 159 407 165 408
rect 31 402 37 403
rect 31 398 32 402
rect 36 398 37 402
rect 31 397 37 398
rect 95 382 101 383
rect 95 378 96 382
rect 100 378 101 382
rect 95 377 101 378
rect 87 372 93 373
rect 87 368 88 372
rect 92 368 93 372
rect 96 369 100 377
rect 87 367 93 368
rect 8 363 12 367
rect 112 361 116 407
rect 119 402 125 403
rect 119 398 120 402
rect 124 398 125 402
rect 119 397 125 398
rect 120 392 125 397
rect 144 378 148 407
rect 151 402 157 403
rect 151 398 152 402
rect 156 398 157 402
rect 151 397 157 398
rect 128 363 132 371
rect 127 362 133 363
rect 127 358 128 362
rect 132 358 133 362
rect 127 357 133 358
rect 152 353 156 397
rect 160 363 164 407
rect 167 372 173 373
rect 167 368 168 372
rect 172 368 173 372
rect 167 367 173 368
rect 15 342 21 343
rect 15 338 16 342
rect 20 338 21 342
rect 15 337 21 338
rect 0 233 4 266
rect 16 247 20 337
rect 111 302 117 303
rect 111 298 112 302
rect 116 298 117 302
rect 111 297 117 298
rect 143 302 149 303
rect 143 298 144 302
rect 148 298 149 302
rect 143 297 149 298
rect 159 302 165 303
rect 159 298 160 302
rect 164 298 165 302
rect 159 297 165 298
rect 31 292 37 293
rect 31 288 32 292
rect 36 288 37 292
rect 95 272 101 273
rect 95 268 96 272
rect 100 268 101 272
rect 95 267 101 268
rect 87 262 93 263
rect 87 258 88 262
rect 92 258 93 262
rect 96 259 100 267
rect 87 257 93 258
rect 112 251 116 297
rect 119 292 125 293
rect 119 288 120 292
rect 124 288 125 292
rect 119 287 125 288
rect 120 285 125 287
rect 120 282 124 285
rect 144 268 148 297
rect 151 292 157 293
rect 151 288 152 292
rect 156 288 157 292
rect 151 287 157 288
rect 128 253 132 261
rect 127 252 133 253
rect 127 248 128 252
rect 132 248 133 252
rect 127 247 133 248
rect 152 243 156 287
rect 160 253 164 297
rect 167 262 173 263
rect 167 258 168 262
rect 172 258 173 262
rect 167 257 173 258
rect -1 232 5 233
rect -1 228 0 232
rect 4 228 5 232
rect -1 227 5 228
rect 111 192 117 193
rect 111 188 112 192
rect 116 188 117 192
rect 111 187 117 188
rect 143 192 149 193
rect 143 188 144 192
rect 148 188 149 192
rect 143 187 149 188
rect 159 192 165 193
rect 159 188 160 192
rect 164 188 165 192
rect 159 187 165 188
rect 95 162 101 163
rect 95 158 96 162
rect 100 158 101 162
rect 95 157 101 158
rect 87 152 93 153
rect 87 148 88 152
rect 92 148 93 152
rect 96 149 100 157
rect 87 147 93 148
rect 112 141 116 187
rect 119 182 125 183
rect 119 178 120 182
rect 124 178 125 182
rect 119 177 125 178
rect 120 175 125 177
rect 120 172 124 175
rect 144 158 148 187
rect 151 182 157 183
rect 151 178 152 182
rect 156 178 157 182
rect 151 177 157 178
rect 128 143 132 151
rect 127 142 133 143
rect 127 138 128 142
rect 132 138 133 142
rect 127 137 133 138
rect 152 133 156 177
rect 160 143 164 187
rect 167 152 173 153
rect 167 148 168 152
rect 172 148 173 152
rect 167 147 173 148
rect 15 122 21 123
rect 15 118 16 122
rect 20 118 21 122
rect 15 117 21 118
rect 0 13 4 46
rect 16 27 20 117
rect 111 82 117 83
rect 111 78 112 82
rect 116 78 117 82
rect 111 77 117 78
rect 143 82 149 83
rect 143 78 144 82
rect 148 78 149 82
rect 143 77 149 78
rect 159 82 165 83
rect 159 78 160 82
rect 164 78 165 82
rect 159 77 165 78
rect 31 72 37 73
rect 31 68 32 72
rect 36 68 37 72
rect 31 67 37 68
rect 95 52 101 53
rect 95 48 96 52
rect 100 48 101 52
rect 95 47 101 48
rect 87 42 93 43
rect 87 38 88 42
rect 92 38 93 42
rect 96 39 100 47
rect 87 37 93 38
rect 112 31 116 77
rect 119 72 125 73
rect 119 68 120 72
rect 124 68 125 72
rect 119 67 125 68
rect 120 65 125 67
rect 120 62 124 65
rect 144 48 148 77
rect 151 72 157 73
rect 151 68 152 72
rect 156 68 157 72
rect 151 67 157 68
rect 128 33 132 41
rect 127 32 133 33
rect 127 28 128 32
rect 132 28 133 32
rect 127 27 133 28
rect 152 23 156 67
rect 160 33 164 77
rect 167 42 173 43
rect 167 38 168 42
rect 172 38 173 42
rect 167 37 173 38
rect 176 23 180 50
rect 192 23 196 917
rect 263 852 269 853
rect 263 848 264 852
rect 268 848 269 852
rect 263 847 269 848
rect 343 852 349 853
rect 343 848 344 852
rect 348 848 349 852
rect 343 847 349 848
rect 264 782 268 847
rect 303 822 309 823
rect 303 818 304 822
rect 308 818 309 822
rect 303 817 309 818
rect 304 805 308 817
rect 344 807 348 847
rect 312 803 316 807
rect 311 802 317 803
rect 311 798 312 802
rect 316 798 317 802
rect 311 797 317 798
rect 263 742 269 743
rect 263 738 264 742
rect 268 738 269 742
rect 263 737 269 738
rect 343 742 349 743
rect 343 738 344 742
rect 348 738 349 742
rect 343 737 349 738
rect 264 672 268 737
rect 303 712 309 713
rect 303 708 304 712
rect 308 708 309 712
rect 344 710 348 737
rect 303 707 309 708
rect 304 695 308 707
rect 312 693 316 697
rect 311 692 317 693
rect 311 688 312 692
rect 316 688 317 692
rect 311 687 317 688
rect 263 632 269 633
rect 263 628 264 632
rect 268 628 269 632
rect 263 627 269 628
rect 343 632 349 633
rect 343 628 344 632
rect 348 628 349 632
rect 343 627 349 628
rect 264 562 268 627
rect 303 602 309 603
rect 303 598 304 602
rect 308 598 309 602
rect 344 600 348 627
rect 303 597 309 598
rect 304 585 308 597
rect 312 583 316 587
rect 311 582 317 583
rect 311 578 312 582
rect 316 578 317 582
rect 311 577 317 578
rect 263 522 269 523
rect 263 518 264 522
rect 268 518 269 522
rect 263 517 269 518
rect 343 522 349 523
rect 343 518 344 522
rect 348 518 349 522
rect 343 517 349 518
rect 264 452 268 517
rect 303 492 309 493
rect 303 488 304 492
rect 308 488 309 492
rect 344 490 348 517
rect 303 487 309 488
rect 304 475 308 487
rect 312 473 316 477
rect 311 472 317 473
rect 311 468 312 472
rect 316 468 317 472
rect 311 467 317 468
rect 263 412 269 413
rect 263 408 264 412
rect 268 408 269 412
rect 263 407 269 408
rect 343 412 349 413
rect 343 408 344 412
rect 348 408 349 412
rect 343 407 349 408
rect 264 342 268 407
rect 303 382 309 383
rect 303 378 304 382
rect 308 378 309 382
rect 344 380 348 407
rect 303 377 309 378
rect 304 365 308 377
rect 312 363 316 367
rect 311 362 317 363
rect 311 358 312 362
rect 316 358 317 362
rect 311 357 317 358
rect 263 302 269 303
rect 263 298 264 302
rect 268 298 269 302
rect 263 297 269 298
rect 343 302 349 303
rect 343 298 344 302
rect 348 298 349 302
rect 343 297 349 298
rect 264 232 268 297
rect 303 272 309 273
rect 303 268 304 272
rect 308 268 309 272
rect 344 270 348 297
rect 303 267 309 268
rect 304 255 308 267
rect 312 253 316 257
rect 311 252 317 253
rect 311 248 312 252
rect 316 248 317 252
rect 311 247 317 248
rect 263 192 269 193
rect 263 188 264 192
rect 268 188 269 192
rect 263 187 269 188
rect 343 192 349 193
rect 343 188 344 192
rect 348 188 349 192
rect 343 187 349 188
rect 264 122 268 187
rect 303 162 309 163
rect 303 158 304 162
rect 308 158 309 162
rect 344 160 348 187
rect 303 157 309 158
rect 304 145 308 157
rect 312 143 316 147
rect 311 142 317 143
rect 311 138 312 142
rect 316 138 317 142
rect 311 137 317 138
rect 263 82 269 83
rect 263 78 264 82
rect 268 78 269 82
rect 263 77 269 78
rect 343 82 349 83
rect 343 78 344 82
rect 348 78 349 82
rect 343 77 349 78
rect 175 22 181 23
rect 175 18 176 22
rect 180 18 181 22
rect 175 17 181 18
rect 191 22 197 23
rect 191 18 192 22
rect 196 18 197 22
rect 191 17 197 18
rect -1 12 5 13
rect 264 12 268 77
rect 303 52 309 53
rect 303 48 304 52
rect 308 48 309 52
rect 344 50 348 77
rect 303 47 309 48
rect 304 35 308 47
rect 352 37 356 803
rect 360 772 364 806
rect 384 783 388 810
rect 383 782 389 783
rect 383 778 384 782
rect 388 778 389 782
rect 383 777 389 778
rect 360 662 364 696
rect 384 673 388 700
rect 383 672 389 673
rect 383 668 384 672
rect 388 668 389 672
rect 383 667 389 668
rect 360 552 364 586
rect 384 563 388 590
rect 383 562 389 563
rect 383 558 384 562
rect 388 558 389 562
rect 383 557 389 558
rect 360 442 364 476
rect 384 453 388 480
rect 383 452 389 453
rect 383 448 384 452
rect 388 448 389 452
rect 383 447 389 448
rect 360 332 364 366
rect 384 343 388 370
rect 383 342 389 343
rect 383 338 384 342
rect 388 338 389 342
rect 383 337 389 338
rect 360 222 364 256
rect 384 233 388 260
rect 383 232 389 233
rect 383 228 384 232
rect 388 228 389 232
rect 383 227 389 228
rect 360 112 364 146
rect 384 123 388 150
rect 383 122 389 123
rect 383 118 384 122
rect 388 118 389 122
rect 383 117 389 118
rect 312 33 316 37
rect 311 32 317 33
rect 311 28 312 32
rect 316 28 317 32
rect 311 27 317 28
rect 384 13 388 40
rect 383 12 389 13
rect -1 8 0 12
rect 4 8 5 12
rect -1 7 5 8
rect 383 8 384 12
rect 388 8 389 12
rect 383 7 389 8
<< m3contact >>
rect 48 918 52 922
rect 192 918 196 922
rect 112 848 116 852
rect 144 848 148 852
rect 160 848 164 852
rect 32 838 36 842
rect 96 818 100 822
rect 88 808 92 812
rect 120 838 124 842
rect 152 838 156 842
rect 128 798 132 802
rect 168 808 172 812
rect 16 778 20 782
rect 112 738 116 742
rect 144 738 148 742
rect 160 738 164 742
rect 32 728 36 732
rect 96 708 100 712
rect 88 698 92 702
rect 120 728 124 732
rect 152 728 156 732
rect 128 688 132 692
rect 168 698 172 702
rect 0 668 4 672
rect 112 628 116 632
rect 144 628 148 632
rect 160 628 164 632
rect 32 618 36 622
rect 96 598 100 602
rect 88 588 92 592
rect 120 618 124 622
rect 152 618 156 622
rect 128 578 132 582
rect 168 588 172 592
rect 0 558 4 562
rect 112 518 116 522
rect 144 518 148 522
rect 160 518 164 522
rect 32 508 36 512
rect 96 488 100 492
rect 88 478 92 482
rect 120 508 124 512
rect 152 508 156 512
rect 128 468 132 472
rect 168 478 172 482
rect 16 448 20 452
rect 112 408 116 412
rect 144 408 148 412
rect 160 408 164 412
rect 32 398 36 402
rect 96 378 100 382
rect 88 368 92 372
rect 120 398 124 402
rect 152 398 156 402
rect 128 358 132 362
rect 168 368 172 372
rect 16 338 20 342
rect 112 298 116 302
rect 144 298 148 302
rect 160 298 164 302
rect 32 288 36 292
rect 96 268 100 272
rect 88 258 92 262
rect 120 288 124 292
rect 152 288 156 292
rect 128 248 132 252
rect 168 258 172 262
rect 0 228 4 232
rect 112 188 116 192
rect 144 188 148 192
rect 160 188 164 192
rect 96 158 100 162
rect 88 148 92 152
rect 120 178 124 182
rect 152 178 156 182
rect 128 138 132 142
rect 168 148 172 152
rect 16 118 20 122
rect 112 78 116 82
rect 144 78 148 82
rect 160 78 164 82
rect 32 68 36 72
rect 96 48 100 52
rect 88 38 92 42
rect 120 68 124 72
rect 152 68 156 72
rect 128 28 132 32
rect 168 38 172 42
rect 264 848 268 852
rect 344 848 348 852
rect 304 818 308 822
rect 312 798 316 802
rect 264 738 268 742
rect 344 738 348 742
rect 304 708 308 712
rect 312 688 316 692
rect 264 628 268 632
rect 344 628 348 632
rect 304 598 308 602
rect 312 578 316 582
rect 264 518 268 522
rect 344 518 348 522
rect 304 488 308 492
rect 312 468 316 472
rect 264 408 268 412
rect 344 408 348 412
rect 304 378 308 382
rect 312 358 316 362
rect 264 298 268 302
rect 344 298 348 302
rect 304 268 308 272
rect 312 248 316 252
rect 264 188 268 192
rect 344 188 348 192
rect 304 158 308 162
rect 312 138 316 142
rect 264 78 268 82
rect 344 78 348 82
rect 176 18 180 22
rect 192 18 196 22
rect 304 48 308 52
rect 384 778 388 782
rect 384 668 388 672
rect 384 558 388 562
rect 384 448 388 452
rect 384 338 388 342
rect 384 228 388 232
rect 384 118 388 122
rect 312 28 316 32
rect 0 8 4 12
rect 384 8 388 12
<< metal3 >>
rect 47 922 197 923
rect 47 918 48 922
rect 52 918 192 922
rect 196 918 197 922
rect 47 917 197 918
rect -17 852 165 853
rect -17 848 112 852
rect 116 848 144 852
rect 148 848 160 852
rect 164 848 165 852
rect -17 847 165 848
rect 263 852 349 853
rect 263 848 264 852
rect 268 848 344 852
rect 348 848 349 852
rect 263 847 349 848
rect -17 842 157 843
rect -17 838 32 842
rect 36 838 120 842
rect 124 838 152 842
rect 156 838 157 842
rect -17 837 157 838
rect 95 822 309 823
rect 95 818 96 822
rect 100 818 304 822
rect 308 818 309 822
rect 95 817 309 818
rect 87 812 173 813
rect 87 808 88 812
rect 92 808 168 812
rect 172 808 173 812
rect 87 807 173 808
rect 127 802 317 803
rect 127 798 128 802
rect 132 798 312 802
rect 316 798 317 802
rect 127 797 317 798
rect -17 782 389 783
rect -17 778 16 782
rect 20 778 384 782
rect 388 778 389 782
rect -17 777 389 778
rect -17 742 165 743
rect -17 738 112 742
rect 116 738 144 742
rect 148 738 160 742
rect 164 738 165 742
rect -17 737 165 738
rect 263 742 349 743
rect 263 738 264 742
rect 268 738 344 742
rect 348 738 349 742
rect 263 737 349 738
rect -17 732 157 733
rect -17 728 32 732
rect 36 728 120 732
rect 124 728 152 732
rect 156 728 157 732
rect -17 727 157 728
rect 95 712 309 713
rect 95 708 96 712
rect 100 708 304 712
rect 308 708 309 712
rect 95 707 309 708
rect 87 702 173 703
rect 87 698 88 702
rect 92 698 168 702
rect 172 698 173 702
rect 87 697 173 698
rect 127 692 317 693
rect 127 688 128 692
rect 132 688 312 692
rect 316 688 317 692
rect 127 687 317 688
rect -17 672 389 673
rect -17 668 0 672
rect 4 668 384 672
rect 388 668 389 672
rect -17 667 389 668
rect -17 632 165 633
rect -17 628 112 632
rect 116 628 144 632
rect 148 628 160 632
rect 164 628 165 632
rect -17 627 165 628
rect 263 632 349 633
rect 263 628 264 632
rect 268 628 344 632
rect 348 628 349 632
rect 263 627 349 628
rect -17 622 157 623
rect -17 618 32 622
rect 36 618 120 622
rect 124 618 152 622
rect 156 618 157 622
rect -17 617 157 618
rect 95 602 309 603
rect 95 598 96 602
rect 100 598 304 602
rect 308 598 309 602
rect 95 597 309 598
rect 87 592 173 593
rect 87 588 88 592
rect 92 588 168 592
rect 172 588 173 592
rect 87 587 173 588
rect 127 582 317 583
rect 127 578 128 582
rect 132 578 312 582
rect 316 578 317 582
rect 127 577 317 578
rect -17 562 389 563
rect -17 558 0 562
rect 4 558 384 562
rect 388 558 389 562
rect -17 557 389 558
rect -17 522 165 523
rect -17 518 112 522
rect 116 518 144 522
rect 148 518 160 522
rect 164 518 165 522
rect -17 517 165 518
rect 263 522 349 523
rect 263 518 264 522
rect 268 518 344 522
rect 348 518 349 522
rect 263 517 349 518
rect -17 512 157 513
rect -17 508 32 512
rect 36 508 120 512
rect 124 508 152 512
rect 156 508 157 512
rect -17 507 157 508
rect 95 492 309 493
rect 95 488 96 492
rect 100 488 304 492
rect 308 488 309 492
rect 95 487 309 488
rect 87 482 173 483
rect 87 478 88 482
rect 92 478 168 482
rect 172 478 173 482
rect 87 477 173 478
rect 127 472 317 473
rect 127 468 128 472
rect 132 468 312 472
rect 316 468 317 472
rect 127 467 317 468
rect -17 452 389 453
rect -17 448 16 452
rect 20 448 384 452
rect 388 448 389 452
rect -17 447 389 448
rect -17 412 165 413
rect -17 408 112 412
rect 116 408 144 412
rect 148 408 160 412
rect 164 408 165 412
rect -17 407 165 408
rect 263 412 349 413
rect 263 408 264 412
rect 268 408 344 412
rect 348 408 349 412
rect 263 407 349 408
rect -17 402 157 403
rect -17 398 32 402
rect 36 398 120 402
rect 124 398 152 402
rect 156 398 157 402
rect -17 397 157 398
rect 95 382 309 383
rect 95 378 96 382
rect 100 378 304 382
rect 308 378 309 382
rect 95 377 309 378
rect 87 372 173 373
rect 87 368 88 372
rect 92 368 168 372
rect 172 368 173 372
rect 87 367 173 368
rect 127 362 317 363
rect 127 358 128 362
rect 132 358 312 362
rect 316 358 317 362
rect 127 357 317 358
rect -17 342 389 343
rect -17 338 16 342
rect 20 338 384 342
rect 388 338 389 342
rect -17 337 389 338
rect -17 302 165 303
rect -17 298 112 302
rect 116 298 144 302
rect 148 298 160 302
rect 164 298 165 302
rect -17 297 165 298
rect 263 302 349 303
rect 263 298 264 302
rect 268 298 344 302
rect 348 298 349 302
rect 263 297 349 298
rect -17 292 157 293
rect -17 288 32 292
rect 36 288 120 292
rect 124 288 152 292
rect 156 288 157 292
rect -17 287 21 288
rect 85 287 157 288
rect 95 272 309 273
rect 95 268 96 272
rect 100 268 304 272
rect 308 268 309 272
rect 95 267 309 268
rect 87 262 173 263
rect 87 258 88 262
rect 92 258 168 262
rect 172 258 173 262
rect 87 257 173 258
rect 127 252 317 253
rect 127 248 128 252
rect 132 248 312 252
rect 316 248 317 252
rect 127 247 317 248
rect -17 232 389 233
rect -17 228 0 232
rect 4 228 384 232
rect 388 228 389 232
rect -17 227 389 228
rect -17 192 165 193
rect -17 188 112 192
rect 116 188 144 192
rect 148 188 160 192
rect 164 188 165 192
rect -17 187 165 188
rect 263 192 349 193
rect 263 188 264 192
rect 268 188 344 192
rect 348 188 349 192
rect 263 187 349 188
rect -17 182 157 183
rect -17 178 120 182
rect 124 178 152 182
rect 156 178 157 182
rect -17 177 157 178
rect 95 162 309 163
rect 95 158 96 162
rect 100 158 304 162
rect 308 158 309 162
rect 95 157 309 158
rect 87 152 173 153
rect 87 148 88 152
rect 92 148 168 152
rect 172 148 173 152
rect 87 147 173 148
rect 127 142 317 143
rect 127 138 128 142
rect 132 138 312 142
rect 316 138 317 142
rect 127 137 317 138
rect -17 122 389 123
rect -17 118 16 122
rect 20 118 384 122
rect 388 118 389 122
rect -17 117 389 118
rect -17 82 165 83
rect -17 78 112 82
rect 116 78 144 82
rect 148 78 160 82
rect 164 78 165 82
rect -17 77 165 78
rect 263 82 349 83
rect 263 78 264 82
rect 268 78 344 82
rect 348 78 349 82
rect 263 77 349 78
rect -17 72 157 73
rect -17 68 32 72
rect 36 68 120 72
rect 124 68 152 72
rect 156 68 157 72
rect -17 67 157 68
rect 95 52 309 53
rect 95 48 96 52
rect 100 48 304 52
rect 308 48 309 52
rect 95 47 309 48
rect 87 42 173 43
rect 87 38 88 42
rect 92 38 168 42
rect 172 38 173 42
rect 87 37 173 38
rect 127 32 317 33
rect 127 28 128 32
rect 132 28 312 32
rect 316 28 317 32
rect 127 27 317 28
rect 175 22 197 23
rect 175 18 176 22
rect 180 18 192 22
rect 196 18 197 22
rect 175 17 197 18
rect -17 12 389 13
rect -17 8 0 12
rect 4 8 384 12
rect 388 8 389 12
rect -17 7 389 8
use yzdetect_8  yzdetect_8_0
timestamp 1484534894
transform 1 0 0 0 1 0
box -8 -4 28 756
use condinv  condinv_0
timestamp 1484534894
transform 1 0 32 0 1 0
box -6 -4 66 976
use or2_1x_8  or2_1x_8_0
timestamp 1484433330
transform 1 0 128 0 1 0
box -6 -4 34 866
use adder_8  adder_8_0
timestamp 1484427118
transform 1 0 160 0 1 0
box -6 -4 130 866
use mux4_1x_8  mux4_1x_8_0
timestamp 1484532969
transform 1 0 288 0 1 0
box -6 -4 106 976
<< labels >>
rlabel metal3 -15 10 -15 10 3 result_0_
rlabel metal3 -15 69 -15 69 3 b_0_
rlabel metal3 -14 80 -14 80 3 a_0_
rlabel metal3 -14 120 -14 120 3 result_1_
rlabel metal3 -14 180 -14 180 3 b_1_
rlabel metal3 -14 190 -14 190 3 a_1_
rlabel metal3 -14 230 -14 230 3 result_2_
rlabel metal3 -14 290 -14 290 3 b_2_
rlabel metal3 -13 300 -13 300 3 a_2_
rlabel metal3 -13 399 -13 399 3 b_3_
rlabel metal3 -15 510 -15 510 3 b_4_
rlabel metal3 -14 520 -14 520 3 a_4_
rlabel metal3 -14 560 -14 560 3 result_5_
rlabel metal3 -13 620 -13 620 3 b_5_
rlabel metal3 -14 630 -14 630 3 a_5_
rlabel metal3 -14 669 -14 669 3 result_6_
rlabel metal3 -13 730 -13 730 3 b_6_
rlabel metal3 -13 739 -13 739 3 a_6_
rlabel metal3 -14 780 -14 780 3 result_7_
rlabel metal3 -14 839 -14 839 3 b_7_
rlabel metal3 -14 850 -14 850 3 a_7_
rlabel metal3 55 920 55 920 1 alucontrol_2_
rlabel metal1 33 860 33 860 1 Vdd!
rlabel metal1 6 549 6 549 1 Gnd!
rlabel metal1 6 530 6 530 1 Vdd!
rlabel metal1 4 219 4 219 1 Gnd!
rlabel metal1 2 200 2 200 1 Vdd!
rlabel metal1 3 109 3 109 1 Gnd!
rlabel metal1 1 90 1 90 1 Vdd!
rlabel metal1 3 -1 3 -1 1 Gnd!
rlabel metal2 288 918 292 922 1 alucontrol_0_
rlabel metal2 320 918 324 922 1 alucontrol_1_
rlabel metal1 3 310 3 310 1 Vdd!
rlabel metal1 5 330 5 330 1 Gnd!
rlabel metal1 4 419 4 419 1 Vdd!
rlabel metal1 5 440 5 440 1 Gnd!
rlabel metal1 2 640 2 640 1 Vdd!
rlabel metal1 1 659 1 659 1 Gnd!
rlabel metal1 2 749 2 749 1 Vdd!
rlabel metal2 8 363 12 367 1 zero
rlabel metal3 -13 340 -13 340 3 result_3_
rlabel metal3 -14 450 -14 450 3 result_4_
rlabel metal3 -14 410 -14 410 3 a_3_
<< end >>
                                                                                   and2_1x_8.mag                                                                                       0000644 �    Asz0000145 00000000227 13046424132 011145  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1486497882
use and2_1x  and2_1x_0
array 0 0 40 0 7 110
timestamp 1484419738
transform 1 0 6 0 1 4
box -6 -4 34 96
<< end >>
                                                                                                                                                                                                                                                                                                                                                                         and2_1x.mag                                                                                         0000644 �    Asz0000145 00000004020 13045417712 010716  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1484419738
<< nwell >>
rect -6 40 34 96
<< ntransistor >>
rect 5 7 7 14
rect 13 7 15 13
rect 18 7 20 13
<< ptransistor >>
rect 5 73 7 83
rect 13 77 15 83
rect 21 77 23 83
<< ndiffusion >>
rect 0 12 5 14
rect 4 8 5 12
rect 0 7 5 8
rect 7 13 12 14
rect 7 12 13 13
rect 7 8 8 12
rect 12 8 13 12
rect 7 7 13 8
rect 15 7 18 13
rect 20 12 25 13
rect 20 8 21 12
rect 20 7 25 8
<< pdiffusion >>
rect 0 82 5 83
rect 4 73 5 82
rect 7 82 13 83
rect 7 73 8 82
rect 12 77 13 82
rect 15 82 21 83
rect 15 78 16 82
rect 20 78 21 82
rect 15 77 21 78
rect 23 82 28 83
rect 23 78 24 82
rect 23 77 28 78
<< ndcontact >>
rect 0 8 4 12
rect 8 8 12 12
rect 21 8 25 12
<< pdcontact >>
rect 0 73 4 82
rect 8 73 12 82
rect 16 78 20 82
rect 24 78 28 82
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
<< polysilicon >>
rect 5 83 7 85
rect 13 83 15 85
rect 21 83 23 85
rect 5 14 7 73
rect 13 54 15 77
rect 13 52 17 54
rect 15 40 17 52
rect 13 38 17 40
rect 13 34 15 38
rect 13 13 15 30
rect 21 21 23 77
rect 18 19 23 21
rect 18 13 20 19
rect 5 5 7 7
rect 13 5 15 7
rect 18 5 20 7
<< polycontact >>
rect 7 44 11 48
rect 12 30 16 34
rect 23 61 27 65
<< metal1 >>
rect -2 92 30 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 30 92
rect -2 86 30 88
rect 0 82 4 83
rect 8 82 12 86
rect 16 82 20 83
rect 0 42 4 73
rect 16 48 20 78
rect 24 82 28 86
rect 24 77 28 78
rect 11 44 27 48
rect 0 12 4 38
rect 23 19 27 44
rect 21 15 27 19
rect 0 7 4 8
rect 8 12 12 14
rect 8 4 12 8
rect 21 12 25 15
rect 21 7 25 8
rect -2 2 30 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 30 2
rect -2 -4 30 -2
<< m2contact >>
rect 25 61 27 65
rect 27 61 29 65
rect 0 38 4 42
rect 16 30 20 34
<< metal2 >>
rect 24 61 25 65
<< labels >>
rlabel m2contact 2 40 2 40 1 y
rlabel m2contact 18 32 18 32 1 a
rlabel m2contact 27 63 27 63 1 b
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel metal1 -1 0 -1 0 3 Gnd!
<< end >>
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                AND2X2.mag                                                                                          0000644 �    Asz0000145 00000003703 13055352531 010365  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1488311641
<< nwell >>
rect -8 48 40 105
<< ntransistor >>
rect 7 6 9 26
rect 12 6 14 26
rect 20 6 22 26
<< ptransistor >>
rect 7 74 9 94
rect 15 74 17 94
rect 23 54 25 94
<< ndiffusion >>
rect 2 25 7 26
rect 6 6 7 25
rect 9 6 12 26
rect 14 25 20 26
rect 14 6 15 25
rect 19 6 20 25
rect 22 25 27 26
rect 22 6 23 25
<< pdiffusion >>
rect 2 93 7 94
rect 6 74 7 93
rect 9 93 15 94
rect 9 74 10 93
rect 14 74 15 93
rect 17 92 23 94
rect 17 74 18 92
rect 22 58 23 92
rect 18 56 23 58
rect 20 54 23 56
rect 25 93 30 94
rect 25 54 26 93
<< ndcontact >>
rect 2 6 6 25
rect 15 6 19 25
rect 23 6 27 25
<< pdcontact >>
rect 2 74 6 93
rect 10 74 14 93
rect 18 58 22 92
rect 26 54 30 93
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 23 94 25 96
rect 7 73 9 74
rect 5 71 9 73
rect 5 41 7 71
rect 6 37 7 41
rect 15 39 17 74
rect 5 30 7 37
rect 16 37 17 39
rect 5 28 9 30
rect 7 26 9 28
rect 12 26 14 35
rect 23 33 25 54
rect 24 31 25 33
rect 20 26 22 29
rect 7 4 9 6
rect 12 4 14 6
rect 20 4 22 6
<< polycontact >>
rect 2 37 6 41
rect 12 35 16 39
rect 20 29 24 33
<< metal1 >>
rect -2 102 34 103
rect 2 98 14 102
rect 18 98 34 102
rect -2 97 34 98
rect 2 93 6 97
rect 10 93 14 94
rect 11 53 14 74
rect 18 92 22 97
rect 18 56 22 58
rect 26 93 30 94
rect 11 50 23 53
rect 10 43 14 47
rect 2 33 6 37
rect 11 39 14 43
rect 11 36 12 39
rect 20 33 23 50
rect 27 47 30 54
rect 26 43 30 47
rect 9 30 20 32
rect 3 29 20 30
rect 3 27 12 29
rect 3 26 6 27
rect 27 26 30 43
rect 2 25 6 26
rect 23 25 30 26
rect 27 21 30 25
rect 15 3 19 6
rect -2 2 34 3
rect 2 -2 14 2
rect 18 -2 34 2
rect -2 -3 34 -2
<< labels >>
flabel metal1 4 100 4 100 4 FreeSans 26 0 0 0 vdd
flabel metal1 4 0 4 0 4 FreeSans 26 0 0 0 gnd
flabel metal1 4 35 4 35 4 FreeSans 26 0 0 0 A
flabel metal1 12 45 12 45 4 FreeSans 26 0 0 0 B
flabel metal1 28 45 28 45 4 FreeSans 26 0 0 0 Y
<< end >>
                                                             AOI21X1.mag                                                                                         0000644 �    Asz0000145 00000003544 13055352531 010456  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1488311641
<< nwell >>
rect -7 48 39 105
<< ntransistor >>
rect 10 6 12 26
rect 15 6 17 26
rect 23 6 25 16
<< ptransistor >>
rect 7 54 9 94
rect 15 54 17 94
rect 23 54 25 94
<< ndiffusion >>
rect 5 25 10 26
rect 9 6 10 25
rect 12 6 15 26
rect 17 25 22 26
rect 17 6 18 25
rect 22 6 23 16
rect 25 15 30 16
rect 25 6 26 15
<< pdiffusion >>
rect 2 92 7 94
rect 6 58 7 92
rect 2 54 7 58
rect 9 60 10 94
rect 14 60 15 94
rect 9 54 15 60
rect 17 93 23 94
rect 17 54 18 93
rect 22 54 23 93
rect 25 93 30 94
rect 25 54 26 93
<< ndcontact >>
rect 5 6 9 25
rect 18 6 22 25
rect 26 6 30 15
<< pdcontact >>
rect 2 58 6 92
rect 10 60 14 94
rect 18 54 22 93
rect 26 54 30 93
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 23 94 25 96
rect 7 49 9 54
rect 4 29 6 47
rect 15 41 17 54
rect 14 37 17 41
rect 4 27 12 29
rect 10 26 12 27
rect 15 26 17 37
rect 23 16 25 54
rect 10 4 12 6
rect 15 4 17 6
rect 23 4 25 6
<< polycontact >>
rect 6 45 10 49
rect 10 37 14 41
rect 25 19 29 23
<< metal1 >>
rect -2 102 34 103
rect 2 98 14 102
rect 18 98 34 102
rect -2 97 34 98
rect 10 94 14 97
rect 2 92 6 94
rect 18 93 22 94
rect 2 57 6 58
rect 2 54 18 57
rect 26 93 30 94
rect 2 45 6 47
rect 26 47 29 54
rect 2 44 10 45
rect 18 44 30 47
rect 2 43 6 44
rect 10 33 14 37
rect 18 26 21 44
rect 26 43 30 44
rect 5 25 9 26
rect 18 25 22 26
rect 26 23 30 27
rect 26 15 30 16
rect 5 3 9 6
rect 26 3 30 6
rect -2 2 34 3
rect 2 -2 14 2
rect 18 -2 34 2
rect -2 -3 34 -2
<< labels >>
flabel metal1 4 0 4 0 4 FreeSans 26 0 0 0 gnd
flabel metal1 4 100 4 100 4 FreeSans 26 0 0 0 vdd
flabel metal1 4 45 4 45 4 FreeSans 26 0 0 0 A
flabel metal1 12 35 12 35 4 FreeSans 26 0 0 0 B
flabel metal1 28 45 28 45 4 FreeSans 26 0 0 0 Y
flabel metal1 28 25 28 25 4 FreeSans 26 0 0 0 C
<< end >>
                                                                                                                                                            condinv.mag                                                                                         0000644 �    Asz0000145 00000006617 13045420162 011131  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1484534894
<< metal1 >>
rect -2 856 22 864
rect 8 816 19 820
rect 8 809 12 816
rect -2 766 22 774
rect -2 746 22 754
rect 8 706 19 710
rect 8 699 12 706
rect -2 656 22 664
rect -2 636 22 644
rect 8 596 19 600
rect 8 589 12 596
rect -2 546 22 554
rect -2 526 22 534
rect 8 486 19 490
rect 8 479 12 486
rect -2 436 22 444
rect -2 416 22 424
rect 8 376 19 380
rect 8 369 12 376
rect -2 326 22 334
rect -2 306 22 314
rect 8 266 19 270
rect 8 259 12 266
rect -2 216 22 224
rect -2 196 22 204
rect 8 156 19 160
rect 8 149 12 156
rect -2 106 22 114
rect -2 86 22 94
rect 8 46 19 50
rect 8 39 12 46
rect -2 -4 22 4
<< m2contact >>
rect 0 808 4 812
rect 0 698 4 702
rect 0 588 4 592
rect 0 478 4 482
rect 0 368 4 372
rect 0 258 4 262
rect 0 148 4 152
rect 0 38 4 42
<< metal2 >>
rect -1 842 5 843
rect -1 838 0 842
rect 4 838 5 842
rect -1 837 5 838
rect 47 842 53 843
rect 47 838 48 842
rect 52 838 53 842
rect 47 837 53 838
rect 0 812 4 837
rect 48 815 52 837
rect -1 732 5 733
rect -1 728 0 732
rect 4 728 5 732
rect -1 727 5 728
rect 47 732 53 733
rect 47 728 48 732
rect 52 728 53 732
rect 47 727 53 728
rect 0 702 4 727
rect 48 705 52 727
rect -1 622 5 623
rect -1 618 0 622
rect 4 618 5 622
rect -1 617 5 618
rect 47 622 53 623
rect 47 618 48 622
rect 52 618 53 622
rect 47 617 53 618
rect 0 592 4 617
rect 48 595 52 617
rect -1 512 5 513
rect -1 508 0 512
rect 4 508 5 512
rect -1 507 5 508
rect 47 512 53 513
rect 47 508 48 512
rect 52 508 53 512
rect 47 507 53 508
rect 0 482 4 507
rect 48 485 52 507
rect -1 402 5 403
rect -1 398 0 402
rect 4 398 5 402
rect -1 397 5 398
rect 47 402 53 403
rect 47 398 48 402
rect 52 398 53 402
rect 47 397 53 398
rect 0 372 4 397
rect 48 375 52 397
rect -1 292 5 293
rect -1 288 0 292
rect 4 288 5 292
rect -1 287 5 288
rect 47 292 53 293
rect 47 288 48 292
rect 52 288 53 292
rect 47 287 53 288
rect 0 262 4 287
rect 48 265 52 287
rect -1 182 5 183
rect -1 178 0 182
rect 4 178 5 182
rect -1 177 5 178
rect 47 182 53 183
rect 47 178 48 182
rect 52 178 53 182
rect 47 177 53 178
rect 0 152 4 177
rect 48 155 52 177
rect -1 72 5 73
rect -1 68 0 72
rect 4 68 5 72
rect -1 67 5 68
rect 47 72 53 73
rect 47 68 48 72
rect 52 68 53 72
rect 47 67 53 68
rect 0 42 4 67
rect 48 45 52 67
<< m3contact >>
rect 0 838 4 842
rect 48 838 52 842
rect 0 728 4 732
rect 48 728 52 732
rect 0 618 4 622
rect 48 618 52 622
rect 0 508 4 512
rect 48 508 52 512
rect 0 398 4 402
rect 48 398 52 402
rect 0 288 4 292
rect 48 288 52 292
rect 0 178 4 182
rect 48 178 52 182
rect 0 68 4 72
rect 48 68 52 72
<< metal3 >>
rect -1 842 53 843
rect -1 838 0 842
rect 4 838 48 842
rect 52 838 53 842
rect -1 837 53 838
rect -1 732 53 733
rect -1 728 0 732
rect 4 728 48 732
rect 52 728 53 732
rect -1 727 53 728
rect -1 622 53 623
rect -1 618 0 622
rect 4 618 48 622
rect 52 618 53 622
rect -1 617 53 618
rect -1 512 53 513
rect -1 508 0 512
rect 4 508 48 512
rect 52 508 53 512
rect -1 507 53 508
rect -1 402 53 403
rect -1 398 0 402
rect 4 398 48 402
rect 52 398 53 402
rect -1 397 53 398
rect -1 292 53 293
rect -1 288 0 292
rect 4 288 48 292
rect 52 288 53 292
rect -1 287 53 288
rect -1 182 53 183
rect -1 178 0 182
rect 4 178 48 182
rect 52 178 53 182
rect -1 177 53 178
rect -1 72 53 73
rect -1 68 0 72
rect 4 68 48 72
rect 52 68 53 72
rect -1 67 53 68
use inv_1x_8  inv_1x_8_0
timestamp 1484534894
transform 1 0 0 0 1 0
box -6 -4 18 866
use mux2_1x_8  mux2_1x_8_0
timestamp 1484532969
transform 1 0 16 0 1 0
box -6 -4 50 976
<< end >>
                                                                                                                 decoder.mag                                                                                         0000644 �    Asz0000145 00000015777 13055341265 011114  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1488306716
<< metal1 >>
rect 30 225 378 240
rect 55 200 353 215
rect 30 187 378 193
rect 226 138 230 148
rect 274 138 278 148
rect 55 87 353 93
rect 55 65 353 80
rect 30 40 378 55
<< metal2 >>
rect 18 277 45 280
rect 322 277 365 280
rect 18 168 21 277
rect 18 3 21 131
rect 30 40 45 240
rect 55 65 70 215
rect 322 168 325 277
rect 186 137 189 151
rect 106 108 109 134
rect 170 109 173 131
rect 218 115 221 151
rect 234 108 237 134
rect 266 109 269 131
rect 282 3 285 134
rect 306 119 309 131
rect 338 65 353 215
rect 363 40 378 240
rect 18 0 45 3
rect 282 0 365 3
<< metal3 >>
rect 17 167 107 172
rect 182 167 326 172
rect 145 147 222 152
rect 0 137 230 142
rect 273 137 408 142
rect 17 127 310 132
rect 89 117 286 122
rect 105 107 318 112
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_0
timestamp 1488306716
transform 1 0 37 0 1 232
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_1
timestamp 1488306716
transform 1 0 370 0 1 232
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_2
timestamp 1488306716
transform 1 0 62 0 1 207
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_3
timestamp 1488306716
transform 1 0 345 0 1 207
box -7 -7 7 7
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_0
timestamp 1488306716
transform 1 0 37 0 1 190
box -7 -2 7 2
use $$M3_M2  $$M3_M2_0
timestamp 1488306716
transform 1 0 20 0 1 170
box -3 -3 3 3
use $$M3_M2  $$M3_M2_7
timestamp 1488306716
transform 1 0 20 0 1 130
box -3 -3 3 3
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_2
timestamp 1488306716
transform 1 0 62 0 1 90
box -7 -2 7 2
use $$M2_M1  $$M2_M1_0
timestamp 1488306716
transform 1 0 105 0 1 170
box -2 -2 2 2
use $$M3_M2  $$M3_M2_1
timestamp 1488306716
transform 1 0 105 0 1 170
box -3 -3 3 3
use $$M3_M2  $$M3_M2_13
timestamp 1488306716
transform 1 0 92 0 1 120
box -3 -3 3 3
use $$M2_M1  $$M2_M1_11
timestamp 1488306716
transform 1 0 92 0 1 117
box -2 -2 2 2
use FILL  FILL_0
timestamp 1488306716
transform -1 0 88 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_3
timestamp 1488306716
transform 1 0 108 0 1 133
box -2 -2 2 2
use $$M3_M2  $$M3_M2_16
timestamp 1488306716
transform 1 0 108 0 1 110
box -3 -3 3 3
use NOR2X1  NOR2X1_0
timestamp 1488306716
transform 1 0 88 0 1 90
box -8 -3 32 105
use FILL  FILL_1
timestamp 1488306716
transform -1 0 120 0 1 90
box -8 -3 16 105
use FILL  FILL_2
timestamp 1488306716
transform -1 0 128 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_2
timestamp 1488306716
transform 1 0 148 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_4
timestamp 1488306716
transform 1 0 148 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_9
timestamp 1488306716
transform 1 0 140 0 1 121
box -2 -2 2 2
use $$M3_M2  $$M3_M2_14
timestamp 1488306716
transform 1 0 140 0 1 120
box -3 -3 3 3
use FILL  FILL_3
timestamp 1488306716
transform -1 0 136 0 1 90
box -8 -3 16 105
use INVX2  INVX2_0
timestamp 1488306716
transform 1 0 136 0 1 90
box -9 -3 26 105
use FILL  FILL_4
timestamp 1488306716
transform -1 0 160 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_1
timestamp 1488306716
transform 1 0 185 0 1 170
box -2 -2 2 2
use $$M3_M2  $$M3_M2_2
timestamp 1488306716
transform 1 0 185 0 1 170
box -3 -3 3 3
use $$M3_M2  $$M3_M2_10
timestamp 1488306716
transform 1 0 172 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_13
timestamp 1488306716
transform 1 0 172 0 1 111
box -2 -2 2 2
use FILL  FILL_5
timestamp 1488306716
transform -1 0 168 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_5
timestamp 1488306716
transform 1 0 188 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_6
timestamp 1488306716
transform 1 0 188 0 1 139
box -2 -2 2 2
use NOR2X1  NOR2X1_1
timestamp 1488306716
transform 1 0 168 0 1 90
box -8 -3 32 105
use FILL  FILL_6
timestamp 1488306716
transform -1 0 200 0 1 90
box -8 -3 16 105
use FILL  FILL_7
timestamp 1488306716
transform -1 0 208 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_6
timestamp 1488306716
transform 1 0 220 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_4
timestamp 1488306716
transform 1 0 228 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_8
timestamp 1488306716
transform 1 0 228 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_12
timestamp 1488306716
transform 1 0 220 0 1 117
box -2 -2 2 2
use FILL  FILL_8
timestamp 1488306716
transform -1 0 216 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_7
timestamp 1488306716
transform 1 0 236 0 1 133
box -2 -2 2 2
use $$M3_M2  $$M3_M2_17
timestamp 1488306716
transform 1 0 236 0 1 110
box -3 -3 3 3
use NOR2X1  NOR2X1_2
timestamp 1488306716
transform 1 0 216 0 1 90
box -8 -3 32 105
use FILL  FILL_9
timestamp 1488306716
transform -1 0 248 0 1 90
box -8 -3 16 105
use FILL  FILL_10
timestamp 1488306716
transform -1 0 256 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_5
timestamp 1488306716
transform 1 0 276 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_9
timestamp 1488306716
transform 1 0 276 0 1 140
box -3 -3 3 3
use $$M3_M2  $$M3_M2_11
timestamp 1488306716
transform 1 0 268 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_14
timestamp 1488306716
transform 1 0 268 0 1 111
box -2 -2 2 2
use FILL  FILL_11
timestamp 1488306716
transform -1 0 264 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_8
timestamp 1488306716
transform 1 0 284 0 1 133
box -2 -2 2 2
use $$M3_M2  $$M3_M2_15
timestamp 1488306716
transform 1 0 284 0 1 120
box -3 -3 3 3
use NOR2X1  NOR2X1_3
timestamp 1488306716
transform 1 0 264 0 1 90
box -8 -3 32 105
use FILL  FILL_12
timestamp 1488306716
transform -1 0 296 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_3
timestamp 1488306716
transform 1 0 324 0 1 170
box -3 -3 3 3
use $$M3_M2  $$M3_M2_12
timestamp 1488306716
transform 1 0 308 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_10
timestamp 1488306716
transform 1 0 308 0 1 121
box -2 -2 2 2
use FILL  FILL_13
timestamp 1488306716
transform -1 0 304 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_15
timestamp 1488306716
transform 1 0 316 0 1 110
box -2 -2 2 2
use $$M3_M2  $$M3_M2_18
timestamp 1488306716
transform 1 0 316 0 1 110
box -3 -3 3 3
use INVX2  INVX2_1
timestamp 1488306716
transform 1 0 304 0 1 90
box -9 -3 26 105
use FILL  FILL_14
timestamp 1488306716
transform -1 0 328 0 1 90
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_1
timestamp 1488306716
transform 1 0 370 0 1 190
box -7 -2 7 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_3
timestamp 1488306716
transform 1 0 345 0 1 90
box -7 -2 7 2
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_4
timestamp 1488306716
transform 1 0 62 0 1 72
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_5
timestamp 1488306716
transform 1 0 345 0 1 72
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_6
timestamp 1488306716
transform 1 0 37 0 1 47
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_7
timestamp 1488306716
transform 1 0 370 0 1 47
box -7 -7 7 7
<< labels >>
flabel metal3 2 140 2 140 4 FreeSans 26 0 0 0 y3
flabel metal2 364 278 364 278 4 FreeSans 26 0 0 0 y1
flabel metal2 44 278 44 278 4 FreeSans 26 0 0 0 y2
flabel metal3 405 140 405 140 4 FreeSans 26 0 0 0 y0
flabel metal2 364 1 364 1 4 FreeSans 26 0 0 0 a[0]
flabel metal2 44 1 44 1 4 FreeSans 26 0 0 0 a[1]
rlabel metal1 193 46 193 46 1 Vdd!
rlabel metal1 193 73 193 73 1 Gnd!
<< end >>
 FILL.mag                                                                                            0000644 �    Asz0000145 00000000634 13055352531 010215  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1488311641
<< nwell >>
rect -8 48 16 105
<< psubstratepcontact >>
rect -2 -2 2 2
rect 6 -2 10 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 6 98 10 102
<< metal1 >>
rect -2 102 10 103
rect 2 98 6 102
rect -2 97 10 98
rect -2 2 10 3
rect 2 -2 6 2
rect -2 -3 10 -2
<< labels >>
flabel metal1 4 100 4 100 4 FreeSans 26 0 0 0 vdd
flabel metal1 4 0 4 0 4 FreeSans 26 0 0 0 gnd
<< end >>
                                                                                                    fulladder.mag                                                                                       0000644 �    Asz0000145 00000014013 13045420314 011417  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1484419411
<< nwell >>
rect -8 40 128 96
<< ntransistor >>
rect 3 7 5 15
rect 11 7 13 15
rect 19 7 21 15
rect 27 7 29 15
rect 35 7 37 15
rect 43 7 45 15
rect 51 7 53 15
rect 59 7 61 15
rect 67 7 69 15
rect 75 7 77 15
rect 83 7 85 15
rect 91 7 93 15
rect 99 7 101 15
rect 115 7 117 15
<< ptransistor >>
rect 3 65 5 81
rect 11 65 13 81
rect 19 65 21 81
rect 27 65 29 81
rect 35 65 37 81
rect 43 65 45 81
rect 51 65 53 81
rect 59 65 61 81
rect 67 65 69 81
rect 75 65 77 81
rect 83 65 85 81
rect 91 65 93 81
rect 99 65 101 81
rect 115 65 117 81
<< ndiffusion >>
rect 2 7 3 15
rect 5 7 6 15
rect 10 7 11 15
rect 13 7 14 15
rect 18 7 19 15
rect 21 7 22 15
rect 26 7 27 15
rect 29 7 35 15
rect 37 7 38 15
rect 42 7 43 15
rect 45 7 46 15
rect 50 7 51 15
rect 53 7 54 15
rect 58 7 59 15
rect 61 7 62 15
rect 66 7 67 15
rect 69 7 70 15
rect 74 7 75 15
rect 77 7 83 15
rect 85 7 91 15
rect 93 7 94 15
rect 98 7 99 15
rect 101 7 102 15
rect 114 7 115 15
rect 117 7 118 15
<< pdiffusion >>
rect -2 80 3 81
rect 2 66 3 80
rect -2 65 3 66
rect 5 72 6 81
rect 10 72 11 81
rect 5 65 11 72
rect 13 80 19 81
rect 13 66 14 80
rect 18 66 19 80
rect 13 65 19 66
rect 21 80 27 81
rect 21 67 22 80
rect 26 67 27 80
rect 21 65 27 67
rect 29 65 35 81
rect 37 80 43 81
rect 37 66 38 80
rect 42 66 43 80
rect 37 65 43 66
rect 45 80 51 81
rect 45 66 46 80
rect 50 66 51 80
rect 45 65 51 66
rect 53 72 54 81
rect 58 72 59 81
rect 53 65 59 72
rect 61 80 67 81
rect 61 66 62 80
rect 66 66 67 80
rect 61 65 67 66
rect 69 80 75 81
rect 69 67 70 80
rect 74 67 75 80
rect 69 65 75 67
rect 77 65 83 81
rect 85 65 91 81
rect 93 80 99 81
rect 93 66 94 80
rect 98 66 99 80
rect 93 65 99 66
rect 101 80 106 81
rect 101 67 102 80
rect 101 65 106 67
rect 110 80 115 81
rect 114 66 115 80
rect 110 65 115 66
rect 117 80 122 81
rect 117 66 118 80
rect 117 65 122 66
<< ndcontact >>
rect -2 7 2 15
rect 6 7 10 15
rect 14 7 18 15
rect 22 7 26 15
rect 38 7 42 15
rect 46 7 50 15
rect 54 7 58 15
rect 62 7 66 15
rect 70 7 74 15
rect 94 7 98 15
rect 102 7 106 15
rect 110 7 114 15
rect 118 7 122 15
<< pdcontact >>
rect -2 66 2 80
rect 6 72 10 81
rect 14 66 18 80
rect 22 67 26 80
rect 38 66 42 80
rect 46 66 50 80
rect 54 72 58 81
rect 62 66 66 80
rect 70 67 74 80
rect 94 66 98 80
rect 102 67 106 80
rect 110 66 114 80
rect 118 66 122 80
<< psubstratepcontact >>
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
<< nsubstratencontact >>
rect -2 88 2 92
rect 6 88 10 92
rect 14 88 18 92
rect 22 88 26 92
rect 30 88 34 92
rect 38 88 42 92
rect 46 88 50 92
rect 54 88 58 92
rect 62 88 66 92
rect 70 88 74 92
rect 78 88 82 92
rect 86 88 90 92
rect 94 88 98 92
rect 102 88 106 92
rect 110 88 114 92
rect 118 88 122 92
<< polysilicon >>
rect 3 81 5 83
rect 11 81 13 83
rect 19 81 21 83
rect 27 81 29 83
rect 35 81 37 83
rect 43 81 45 83
rect 51 81 53 83
rect 59 81 61 83
rect 67 81 69 83
rect 75 81 77 83
rect 83 81 85 83
rect 91 81 93 83
rect 99 81 101 83
rect 115 81 117 83
rect 3 36 5 65
rect 11 43 13 65
rect 19 51 21 65
rect 3 15 5 32
rect 11 15 13 39
rect 19 15 21 47
rect 27 43 29 65
rect 27 15 29 39
rect 35 36 37 65
rect 43 36 45 65
rect 51 43 53 65
rect 59 51 61 65
rect 35 15 37 32
rect 43 15 45 32
rect 51 15 53 39
rect 59 15 61 47
rect 67 29 69 65
rect 75 51 77 65
rect 67 15 69 25
rect 75 15 77 47
rect 83 43 85 65
rect 83 15 85 39
rect 91 36 93 65
rect 91 15 93 32
rect 99 22 101 65
rect 115 29 117 65
rect 99 15 101 18
rect 115 15 117 25
rect 3 5 5 7
rect 11 5 13 7
rect 19 5 21 7
rect 27 5 29 7
rect 35 5 37 7
rect 43 5 45 7
rect 51 5 53 7
rect 59 5 61 7
rect 67 5 69 7
rect 75 5 77 7
rect 83 5 85 7
rect 91 5 93 7
rect 99 5 101 7
rect 115 5 117 7
<< polycontact >>
rect 18 47 22 51
rect 10 39 14 43
rect 2 32 6 36
rect 26 39 30 43
rect 58 47 62 51
rect 50 39 54 43
rect 34 32 38 36
rect 42 32 46 36
rect 74 47 78 51
rect 66 25 70 29
rect 82 39 86 43
rect 90 32 94 36
rect 114 25 118 29
rect 98 18 102 22
<< metal1 >>
rect -4 92 124 94
rect -4 88 -2 92
rect 2 88 6 92
rect 10 88 14 92
rect 18 88 22 92
rect 26 88 30 92
rect 34 88 38 92
rect 42 88 46 92
rect 50 88 54 92
rect 58 88 62 92
rect 66 88 70 92
rect 74 88 78 92
rect 82 88 86 92
rect 90 88 94 92
rect 98 88 102 92
rect 106 88 110 92
rect 114 88 118 92
rect 122 88 124 92
rect -4 86 124 88
rect 6 81 10 86
rect -2 80 2 81
rect 14 80 18 81
rect 2 66 14 69
rect -2 65 18 66
rect 22 80 26 81
rect 38 80 42 86
rect 54 81 58 86
rect 38 65 42 66
rect 46 80 50 81
rect 62 80 66 81
rect 50 66 62 69
rect 46 65 66 66
rect 70 80 74 81
rect 94 80 98 86
rect 94 65 98 66
rect 102 80 106 81
rect 110 80 114 86
rect 110 65 114 66
rect 118 80 122 81
rect 118 59 122 66
rect 18 55 118 59
rect 22 47 58 51
rect 62 47 74 51
rect 14 39 26 43
rect 30 39 50 43
rect 54 39 82 43
rect 6 32 34 36
rect 38 32 42 36
rect 46 32 90 36
rect 26 25 66 29
rect 70 25 114 29
rect -2 18 18 22
rect -2 15 2 18
rect 14 15 18 18
rect 22 15 26 25
rect 46 18 66 22
rect 46 15 50 18
rect 62 15 66 18
rect 74 18 98 22
rect 70 15 74 18
rect 6 4 10 7
rect 38 4 42 7
rect 54 4 58 7
rect 94 4 98 7
rect 110 4 114 7
rect -4 2 124 4
rect -4 -2 -2 2
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 124 2
rect -4 -4 124 -2
<< m2contact >>
rect 22 67 26 69
rect 22 65 26 67
rect 70 67 74 69
rect 70 65 74 67
rect 102 67 106 69
rect 102 65 106 67
rect 14 55 18 59
rect 118 55 122 59
rect 14 47 18 51
rect 6 39 10 43
rect -2 32 2 36
rect 22 25 26 29
rect 70 18 74 22
rect 102 11 106 15
rect 118 11 122 15
<< metal2 >>
rect 22 29 26 65
rect 70 22 74 65
rect 102 15 106 65
rect 118 15 122 55
<< labels >>
rlabel m2contact 0 34 0 34 1 a
rlabel m2contact 8 41 8 41 1 b
rlabel m2contact 16 49 16 49 1 c
rlabel m2contact 16 57 16 57 1 cout
rlabel m2contact 104 13 104 13 1 s
rlabel metal1 4 89 4 89 1 Vdd!
rlabel metal1 4 -1 4 -1 1 Gnd!
<< end >>
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     inv_1x_8.mag                                                                                        0000644 �    Asz0000145 00000001276 13045422315 011122  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1484534894
use inv_1x  inv_1x_0
timestamp 1484418501
transform 1 0 0 0 1 770
box -6 -4 18 96
use inv_1x  inv_1x_1
timestamp 1484418501
transform 1 0 0 0 1 660
box -6 -4 18 96
use inv_1x  inv_1x_2
timestamp 1484418501
transform 1 0 0 0 1 550
box -6 -4 18 96
use inv_1x  inv_1x_3
timestamp 1484418501
transform 1 0 0 0 1 440
box -6 -4 18 96
use inv_1x  inv_1x_4
timestamp 1484418501
transform 1 0 0 0 1 330
box -6 -4 18 96
use inv_1x  inv_1x_5
timestamp 1484418501
transform 1 0 0 0 1 220
box -6 -4 18 96
use inv_1x  inv_1x_6
timestamp 1484418501
transform 1 0 0 0 1 110
box -6 -4 18 96
use inv_1x  inv_1x_7
timestamp 1484418501
transform 1 0 0 0 1 0
box -6 -4 18 96
<< end >>
                                                                                                                                                                                                                                                                                                                                  inv_1x.mag                                                                                          0000644 �    Asz0000145 00000002113 13045422322 010660  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1484418501
<< nwell >>
rect -6 40 18 96
<< ntransistor >>
rect 5 7 7 14
<< ptransistor >>
rect 5 73 7 83
<< ndiffusion >>
rect 0 12 5 14
rect 4 8 5 12
rect 0 7 5 8
rect 7 12 12 14
rect 7 8 8 12
rect 7 7 12 8
<< pdiffusion >>
rect 0 82 5 83
rect 4 73 5 82
rect 7 82 12 83
rect 7 73 8 82
<< ndcontact >>
rect 0 8 4 12
rect 8 8 12 12
<< pdcontact >>
rect 0 73 4 82
rect 8 73 12 82
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
<< polysilicon >>
rect 5 83 7 85
rect 5 14 7 73
rect 5 5 7 7
<< polycontact >>
rect 1 38 5 42
<< metal1 >>
rect -2 92 14 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 14 92
rect -2 86 14 88
rect 0 82 4 86
rect 8 82 12 83
rect 8 42 12 73
rect 0 12 4 14
rect 0 4 4 8
rect 8 12 12 38
rect 8 7 12 8
rect -2 2 14 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 14 2
rect -2 -4 14 -2
<< m2contact >>
rect 0 38 1 42
rect 1 38 4 42
rect 8 38 12 42
<< labels >>
rlabel m2contact 1 40 1 40 1 a
rlabel m2contact 10 40 10 40 1 y
rlabel metal1 -1 0 -1 0 3 Gnd!
rlabel metal1 -1 90 -1 90 3 Vdd!
<< end >>
                                                                                                                                                                                                                                                                                                                                                                                                                                                     invbuf_4x.mag                                                                                       0000644 �    Asz0000145 00000003532 13045417774 011405  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1484532969
<< nwell >>
rect -6 40 34 96
<< ntransistor >>
rect 5 7 7 34
rect 21 7 23 34
<< ptransistor >>
rect 5 46 7 83
rect 21 46 23 83
<< ndiffusion >>
rect 0 32 5 34
rect 4 8 5 32
rect 0 7 5 8
rect 7 32 12 34
rect 7 8 8 32
rect 7 7 12 8
rect 16 32 21 34
rect 20 8 21 32
rect 16 7 21 8
rect 23 32 28 34
rect 23 8 24 32
rect 23 7 28 8
<< pdiffusion >>
rect 0 81 5 83
rect 4 47 5 81
rect 0 46 5 47
rect 7 81 12 83
rect 7 47 8 81
rect 7 46 12 47
rect 16 81 21 83
rect 20 47 21 81
rect 16 46 21 47
rect 23 81 28 83
rect 23 47 24 81
rect 23 46 28 47
<< ndcontact >>
rect 0 8 4 32
rect 8 8 12 32
rect 16 8 20 32
rect 24 8 28 32
<< pdcontact >>
rect 0 47 4 81
rect 8 47 12 81
rect 16 47 20 81
rect 24 47 28 81
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
<< polysilicon >>
rect 5 83 7 85
rect 21 83 23 85
rect 5 34 7 46
rect 21 41 23 46
rect 17 39 23 41
rect 21 34 23 39
rect 5 5 7 7
rect 21 5 23 7
<< polycontact >>
rect 1 38 5 42
rect 13 38 17 42
<< metal1 >>
rect -2 92 30 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 30 92
rect -2 86 30 88
rect 0 81 4 86
rect 0 46 4 47
rect 8 81 12 83
rect 8 42 12 47
rect 16 81 20 86
rect 16 46 20 47
rect 24 81 28 83
rect 24 42 28 47
rect 12 38 13 42
rect 0 32 4 34
rect 0 4 4 8
rect 8 32 12 38
rect 8 7 12 8
rect 16 32 20 34
rect 16 4 20 8
rect 24 32 28 38
rect 24 7 28 8
rect -2 2 30 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 30 2
rect -2 -4 30 -2
<< m2contact >>
rect 0 38 1 42
rect 1 38 4 42
rect 8 38 12 42
rect 24 38 28 42
<< labels >>
rlabel m2contact 1 40 1 40 1 s
rlabel m2contact 10 40 10 40 1 sb_out
rlabel m2contact 26 40 26 40 1 s_out
rlabel metal1 -1 0 -1 0 3 Gnd!
rlabel metal1 -1 90 -1 90 3 Vdd!
<< end >>
                                                                                                                                                                      INVX2.mag                                                                                           0000644 �    Asz0000145 00000001757 13055352531 010344  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1488311641
<< nwell >>
rect -9 48 26 105
<< ntransistor >>
rect 7 6 9 26
<< ptransistor >>
rect 7 54 9 94
<< ndiffusion >>
rect 2 25 7 26
rect 6 6 7 25
rect 9 25 14 26
rect 9 6 10 25
<< pdiffusion >>
rect 2 93 7 94
rect 6 54 7 93
rect 9 93 14 94
rect 9 54 10 93
<< ndcontact >>
rect 2 6 6 25
rect 10 6 14 25
<< pdcontact >>
rect 2 54 6 93
rect 10 54 14 93
<< psubstratepcontact >>
rect -2 -2 2 2
<< nsubstratencontact >>
rect -2 98 2 102
<< polysilicon >>
rect 7 94 9 96
rect 7 33 9 54
rect 6 29 9 33
rect 7 26 9 29
rect 7 4 9 6
<< polycontact >>
rect 2 29 6 33
<< metal1 >>
rect -2 102 18 103
rect 2 98 18 102
rect -2 97 18 98
rect 2 93 6 97
rect 10 93 14 94
rect 2 33 6 37
rect 2 25 6 26
rect 10 25 14 54
rect 2 3 6 6
rect -2 2 18 3
rect 2 -2 18 2
rect -2 -3 18 -2
<< labels >>
flabel metal1 4 100 4 100 4 FreeSans 26 0 0 0 vdd
flabel metal1 4 0 4 0 4 FreeSans 26 0 0 0 gnd
flabel metal1 12 45 12 45 4 FreeSans 26 0 0 0 Y
flabel metal1 4 35 4 35 4 FreeSans 26 0 0 0 A
<< end >>
                 $$M2_M1_1500_1500_3_1.mag                                                                           0000644 �    Asz0000145 00000000117 13055352531 012162  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1488311641
<< m2contact >>
rect -7 -2 7 2
<< end >>
                                                                                                                                                                                                                                                                                                                                                                                                                                                 $$M2_M1_1500_1500_3_3.mag                                                                           0000644 �    Asz0000145 00000000117 13055352531 012164  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1488311641
<< m2contact >>
rect -7 -7 7 7
<< end >>
                                                                                                                                                                                                                                                                                                                                                                                                                                                 $$M2_M1.mag                                                                                         0000644 �    Asz0000145 00000000117 13055352531 010406  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1488311641
<< m2contact >>
rect -2 -2 2 2
<< end >>
                                                                                                                                                                                                                                                                                                                                                                                                                                                 $$M3_M2.mag                                                                                         0000644 �    Asz0000145 00000000230 13055352531 010404  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1488311641
<< m3contact >>
rect -2 -2 2 2
<< metal3 >>
rect -3 2 3 3
rect -3 -2 -2 2
rect 2 -2 3 2
rect -3 -3 3 -2
<< end >>
                                                                                                                                                                                                                                                                                                                                                                        mux2_1x_8.mag                                                                                       0000644 �    Asz0000145 00000001606 13045417727 011231  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1484532969
<< metal2 >>
rect 8 47 12 921
rect 24 56 28 921
use invbuf_4x  invbuf_4x_0
timestamp 1484532969
transform 1 0 0 0 1 880
box -6 -4 34 96
use mux2_dp_1x  mux2_dp_1x_0
timestamp 1484435125
transform 1 0 0 0 1 770
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_1
timestamp 1484435125
transform 1 0 0 0 1 660
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_2
timestamp 1484435125
transform 1 0 0 0 1 550
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_3
timestamp 1484435125
transform 1 0 0 0 1 440
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_4
timestamp 1484435125
transform 1 0 0 0 1 330
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_5
timestamp 1484435125
transform 1 0 0 0 1 220
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_6
timestamp 1484435125
transform 1 0 0 0 1 110
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_7
timestamp 1484435125
transform 1 0 0 0 1 0
box -6 -4 50 96
<< end >>
                                                                                                                          mux2_dp_1x.mag                                                                                      0000644 �    Asz0000145 00000006015 13045417774 011466  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1484435125
<< nwell >>
rect -6 40 50 96
<< ntransistor >>
rect 10 7 12 13
rect 15 7 17 13
rect 23 7 25 13
rect 28 7 30 13
rect 36 7 38 14
<< ptransistor >>
rect 10 74 12 83
rect 15 74 17 83
rect 23 74 25 83
rect 28 74 30 83
rect 36 73 38 83
<< ndiffusion >>
rect 31 13 36 14
rect 5 12 10 13
rect 9 8 10 12
rect 5 7 10 8
rect 12 7 15 13
rect 17 12 23 13
rect 17 8 18 12
rect 22 8 23 12
rect 17 7 23 8
rect 25 7 28 13
rect 30 12 36 13
rect 30 8 31 12
rect 35 8 36 12
rect 30 7 36 8
rect 38 12 43 14
rect 38 8 39 12
rect 38 7 43 8
<< pdiffusion >>
rect 9 74 10 83
rect 12 74 15 83
rect 17 74 18 83
rect 22 74 23 83
rect 25 74 28 83
rect 30 82 36 83
rect 30 74 31 82
rect 35 73 36 82
rect 38 82 43 83
rect 38 73 39 82
<< ndcontact >>
rect 5 8 9 12
rect 18 8 22 12
rect 31 8 35 12
rect 39 8 43 12
<< pdcontact >>
rect 5 74 9 83
rect 18 74 22 83
rect 31 73 35 82
rect 39 73 43 82
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
rect 40 -2 44 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
rect 32 88 36 92
rect 40 88 44 92
<< polysilicon >>
rect 10 83 12 85
rect 15 83 17 85
rect 23 83 25 85
rect 28 83 30 85
rect 36 83 38 85
rect 10 65 12 74
rect 2 63 12 65
rect 2 50 4 63
rect 15 60 17 74
rect 9 58 17 60
rect 9 50 11 58
rect 23 55 25 74
rect 18 53 25 55
rect 28 49 30 74
rect 2 16 4 46
rect 18 42 20 49
rect 15 40 20 42
rect 2 14 12 16
rect 10 13 12 14
rect 15 13 17 40
rect 27 33 29 45
rect 36 41 38 73
rect 37 37 38 41
rect 27 31 31 33
rect 23 13 25 23
rect 29 17 31 31
rect 28 15 31 17
rect 28 13 30 15
rect 36 14 38 37
rect 10 5 12 7
rect 15 5 17 7
rect 23 5 25 7
rect 28 5 30 7
rect 36 5 38 7
<< polycontact >>
rect 0 46 4 50
rect 8 46 12 50
rect 18 49 22 53
rect 26 45 30 49
rect 33 37 37 41
rect 21 23 25 27
<< metal1 >>
rect -2 92 46 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 32 92
rect 36 88 40 92
rect 44 88 46 92
rect -2 86 46 88
rect 5 83 9 86
rect 18 69 22 74
rect 31 82 35 86
rect 39 82 43 83
rect 20 65 22 69
rect 18 55 24 59
rect 18 53 22 55
rect 39 50 43 73
rect 8 27 12 46
rect 30 45 32 48
rect 26 44 32 45
rect 39 46 44 50
rect 40 42 44 46
rect 31 37 33 41
rect 31 35 35 37
rect 20 32 35 35
rect 20 31 27 32
rect 31 31 35 32
rect 40 31 44 38
rect 39 27 44 31
rect 8 23 21 27
rect 20 15 22 19
rect 5 12 9 13
rect 5 4 9 8
rect 18 12 22 15
rect 18 7 22 8
rect 31 12 35 14
rect 31 4 35 8
rect 39 12 43 27
rect 39 7 43 8
rect -2 2 46 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 40 2
rect 44 -2 46 2
rect -2 -4 46 -2
<< m2contact >>
rect 16 65 20 69
rect 24 55 28 59
rect 0 46 4 50
rect 8 46 12 50
rect 32 44 36 48
rect 40 38 44 42
rect 16 31 20 35
rect 16 15 20 19
<< metal2 >>
rect 16 35 20 65
rect 16 19 20 31
<< labels >>
rlabel metal1 -1 0 -1 0 2 Gnd!
rlabel m2contact 42 40 42 40 1 y
rlabel m2contact 34 46 34 46 1 d0
rlabel m2contact 26 57 26 57 1 s
rlabel m2contact 10 48 10 48 1 sb
rlabel m2contact 2 48 2 48 1 d1
rlabel metal1 -1 90 -1 90 3 Vdd!
<< end >>
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   mux3_1x_8.mag                                                                                       0000644 �    Asz0000145 00000003517 13045677255 011241  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1484532969
<< metal1 >>
rect -2 966 38 974
rect -2 876 38 884
rect 12 868 24 872
rect 44 868 56 872
<< m2contact >>
rect 8 868 12 872
rect 24 868 28 872
rect 40 868 44 872
rect 56 868 60 872
<< metal2 >>
rect -1 902 5 903
rect -1 898 0 902
rect 4 898 5 902
rect -1 897 5 898
rect 0 49 4 897
rect 8 872 12 923
rect 24 903 28 921
rect 40 903 44 921
rect 23 902 29 903
rect 23 898 24 902
rect 28 898 29 902
rect 23 897 29 898
rect 38 902 44 903
rect 38 898 39 902
rect 43 898 44 902
rect 38 897 44 898
rect 47 902 53 903
rect 47 898 48 902
rect 52 898 53 902
rect 47 897 53 898
rect 24 49 28 868
rect 40 40 44 868
rect 48 49 52 897
rect 56 872 60 922
<< m3contact >>
rect 0 898 4 902
rect 24 898 28 902
rect 39 898 43 902
rect 48 898 52 902
<< metal3 >>
rect -1 902 29 903
rect -1 898 0 902
rect 4 898 24 902
rect 28 898 29 902
rect -1 897 29 898
rect 38 902 53 903
rect 38 898 39 902
rect 43 898 48 902
rect 52 898 53 902
rect 38 897 53 898
use invbuf_4x  invbuf_4x_0
timestamp 1484532969
transform 1 0 0 0 1 880
box -6 -4 34 96
use invbuf_4x  invbuf_4x_1
timestamp 1484532969
transform 1 0 32 0 1 880
box -6 -4 34 96
use mux3_dp_1x  mux3_dp_1x_0
timestamp 1484514831
transform 1 0 0 0 1 770
box -6 -4 82 96
use mux3_dp_1x  mux3_dp_1x_1
timestamp 1484514831
transform 1 0 0 0 1 660
box -6 -4 82 96
use mux3_dp_1x  mux3_dp_1x_2
timestamp 1484514831
transform 1 0 0 0 1 550
box -6 -4 82 96
use mux3_dp_1x  mux3_dp_1x_3
timestamp 1484514831
transform 1 0 0 0 1 440
box -6 -4 82 96
use mux3_dp_1x  mux3_dp_1x_4
timestamp 1484514831
transform 1 0 0 0 1 330
box -6 -4 82 96
use mux3_dp_1x  mux3_dp_1x_5
timestamp 1484514831
transform 1 0 0 0 1 220
box -6 -4 82 96
use mux3_dp_1x  mux3_dp_1x_6
timestamp 1484514831
transform 1 0 0 0 1 110
box -6 -4 82 96
use mux3_dp_1x  mux3_dp_1x_7
timestamp 1484514831
transform 1 0 0 0 1 0
box -6 -4 82 96
<< end >>
                                                                                                                                                                                 mux3_dp_1x.mag                                                                                      0000644 �    Asz0000145 00000011226 13045677255 011471  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1484514831
<< nwell >>
rect -6 40 82 96
<< ntransistor >>
rect 5 7 7 13
rect 10 7 12 13
rect 18 7 20 13
rect 23 7 25 13
rect 31 7 33 13
rect 39 7 41 13
rect 44 7 46 13
rect 62 12 69 14
<< ptransistor >>
rect 5 74 7 83
rect 10 74 12 83
rect 18 74 20 83
rect 23 74 25 83
rect 31 74 33 83
rect 39 74 41 83
rect 44 74 46 83
rect 59 73 69 75
<< ndiffusion >>
rect 62 15 63 19
rect 67 15 69 19
rect 62 14 69 15
rect 0 12 5 13
rect 4 8 5 12
rect 0 7 5 8
rect 7 7 10 13
rect 12 12 18 13
rect 12 8 13 12
rect 17 8 18 12
rect 12 7 18 8
rect 20 7 23 13
rect 25 12 31 13
rect 25 8 26 12
rect 30 8 31 12
rect 25 7 31 8
rect 33 12 39 13
rect 33 8 34 12
rect 38 8 39 12
rect 33 7 39 8
rect 41 7 44 13
rect 46 12 51 13
rect 46 8 47 12
rect 46 7 51 8
rect 62 11 69 12
rect 62 7 63 11
rect 67 7 69 11
<< pdiffusion >>
rect 4 74 5 83
rect 7 74 10 83
rect 12 74 13 83
rect 17 74 18 83
rect 20 74 23 83
rect 25 74 26 83
rect 30 74 31 83
rect 33 74 34 83
rect 38 74 39 83
rect 41 74 44 83
rect 46 74 47 83
rect 68 76 69 80
rect 59 75 69 76
rect 59 72 69 73
rect 68 68 69 72
<< ndcontact >>
rect 63 15 67 19
rect 0 8 4 12
rect 13 8 17 12
rect 26 8 30 12
rect 34 8 38 12
rect 47 8 51 12
rect 63 7 67 11
<< pdcontact >>
rect 0 74 4 83
rect 13 74 17 83
rect 26 74 30 83
rect 34 74 38 83
rect 47 74 51 83
rect 59 76 68 80
rect 59 68 68 72
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
rect 40 -2 44 2
rect 48 -2 52 2
rect 56 -2 60 2
rect 64 -2 68 2
rect 72 -2 76 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
rect 32 88 36 92
rect 40 88 44 92
rect 48 88 52 92
rect 56 88 60 92
rect 64 88 68 92
rect 72 88 76 92
<< polysilicon >>
rect 5 83 7 85
rect 10 83 12 85
rect 18 83 20 85
rect 23 83 25 85
rect 31 83 33 85
rect 39 83 41 85
rect 44 83 46 85
rect 5 64 7 74
rect 0 62 7 64
rect 0 52 2 62
rect 10 58 12 74
rect 18 64 20 74
rect 9 56 12 58
rect 16 62 20 64
rect 0 26 2 48
rect 9 43 11 56
rect 16 52 18 62
rect 23 59 25 74
rect 31 73 33 74
rect 31 71 36 73
rect 23 57 30 59
rect 28 49 30 57
rect 34 54 36 71
rect 39 59 41 74
rect 44 64 46 74
rect 57 73 59 75
rect 69 73 72 75
rect 44 62 59 64
rect 70 62 72 73
rect 39 57 50 59
rect 34 52 42 54
rect 16 32 18 48
rect 28 47 35 49
rect 23 32 25 39
rect 33 35 35 47
rect 40 43 42 52
rect 48 52 50 57
rect 57 52 59 62
rect 67 58 72 62
rect 60 48 65 51
rect 13 30 18 32
rect 21 30 25 32
rect 29 33 35 35
rect 48 34 50 48
rect 0 24 7 26
rect 5 13 7 24
rect 13 16 15 30
rect 21 27 23 30
rect 29 27 31 33
rect 44 32 50 34
rect 44 30 46 32
rect 10 14 15 16
rect 18 25 23 27
rect 26 25 31 27
rect 34 28 46 30
rect 55 28 57 39
rect 10 13 12 14
rect 18 13 20 25
rect 26 16 28 25
rect 34 22 36 28
rect 53 26 57 28
rect 53 25 55 26
rect 23 14 28 16
rect 31 20 36 22
rect 39 23 55 25
rect 23 13 25 14
rect 31 13 33 20
rect 39 13 41 23
rect 63 22 65 48
rect 59 20 65 22
rect 44 18 61 20
rect 44 13 46 18
rect 70 14 72 58
rect 60 12 62 14
rect 69 12 72 14
rect 5 5 7 7
rect 10 5 12 7
rect 18 5 20 7
rect 23 5 25 7
rect 31 5 33 7
rect 39 5 41 7
rect 44 5 46 7
<< polycontact >>
rect 0 48 4 52
rect 16 48 20 52
rect 24 48 28 52
rect 8 39 12 43
rect 22 39 26 43
rect 63 58 67 62
rect 48 48 52 52
rect 56 48 60 52
rect 40 39 44 43
rect 54 39 58 43
<< metal1 >>
rect -2 92 78 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 32 92
rect 36 88 40 92
rect 44 88 48 92
rect 52 88 56 92
rect 60 88 64 92
rect 68 88 72 92
rect 76 88 78 92
rect -2 86 78 88
rect 13 83 17 86
rect 47 83 51 86
rect 0 70 4 74
rect 26 70 30 74
rect 0 66 30 70
rect 62 80 66 86
rect 68 76 69 80
rect 0 58 4 66
rect 34 62 38 74
rect 68 68 76 72
rect 34 58 63 62
rect 12 39 22 43
rect 44 39 54 43
rect 63 28 67 58
rect 34 24 67 28
rect 72 42 76 68
rect 0 17 30 21
rect 0 12 4 17
rect 0 7 4 8
rect 13 12 17 13
rect 13 4 17 8
rect 26 12 30 17
rect 26 7 30 8
rect 34 12 38 24
rect 72 19 76 38
rect 62 15 63 19
rect 67 15 76 19
rect 34 7 38 8
rect 47 12 51 13
rect 47 4 51 8
rect 62 7 63 11
rect 67 7 69 11
rect 63 4 67 7
rect -2 2 78 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 40 2
rect 44 -2 48 2
rect 52 -2 56 2
rect 60 -2 64 2
rect 68 -2 72 2
rect 76 -2 78 2
rect -2 -4 78 -2
<< m2contact >>
rect 0 48 4 52
rect 16 48 20 52
rect 24 48 28 52
rect 48 48 52 52
rect 56 48 60 52
rect 8 39 12 43
rect 40 39 44 43
rect 72 38 76 42
<< labels >>
rlabel m2contact 2 50 2 50 1 s0
rlabel m2contact 18 50 18 50 1 d1
rlabel m2contact 26 50 26 50 1 s0b
rlabel m2contact 50 50 50 50 1 s1b
rlabel m2contact 58 50 58 50 1 d2
rlabel m2contact 74 40 74 40 1 y
rlabel m2contact 42 41 42 41 1 s1
rlabel m2contact 10 41 10 41 1 d0
rlabel metal1 -1 89 -1 89 3 Vdd!
rlabel metal1 -1 0 -1 0 2 Gnd!
<< end >>
                                                                                                                                                                                                                                                                                                                                                                          mux4_1x_8.mag                                                                                       0000644 �    Asz0000145 00000004232 13045420406 011215  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1484532969
<< metal1 >>
rect -2 966 38 974
rect -2 876 38 884
rect 4 868 8 872
rect 44 868 48 872
<< m2contact >>
rect 0 868 4 872
rect 8 868 12 872
rect 40 868 44 872
rect 48 868 52 872
<< metal2 >>
rect 0 918 4 922
rect 8 872 12 922
rect 24 913 28 921
rect 32 918 36 922
rect 23 912 29 913
rect 23 908 24 912
rect 28 908 29 912
rect 23 907 29 908
rect 31 902 37 903
rect 31 898 32 902
rect 36 898 37 902
rect 31 897 37 898
rect 0 43 4 868
rect 32 50 36 897
rect 40 872 44 922
rect 56 903 60 921
rect 79 912 85 913
rect 79 908 80 912
rect 84 908 85 912
rect 79 907 85 908
rect 55 902 61 903
rect 55 898 56 902
rect 60 898 61 902
rect 55 897 61 898
rect 16 34 20 38
rect 24 34 28 38
rect 48 35 52 868
rect 80 57 84 907
rect 96 37 100 41
rect 72 33 76 37
<< m3contact >>
rect 24 908 28 912
rect 32 898 36 902
rect 80 908 84 912
rect 56 898 60 902
<< metal3 >>
rect 23 912 85 913
rect 23 908 24 912
rect 28 908 80 912
rect 84 908 85 912
rect 23 907 85 908
rect 31 902 61 903
rect 31 898 32 902
rect 36 898 56 902
rect 60 898 61 902
rect 31 897 61 898
use invbuf_4x  invbuf_4x_0
timestamp 1484532969
transform 1 0 0 0 1 880
box -6 -4 34 96
use invbuf_4x  invbuf_4x_1
timestamp 1484532969
transform 1 0 32 0 1 880
box -6 -4 34 96
use mux4_dp_1x  mux4_dp_1x_0
timestamp 1484419186
transform 1 0 0 0 1 770
box -6 -4 106 96
use mux4_dp_1x  mux4_dp_1x_1
timestamp 1484419186
transform 1 0 0 0 1 660
box -6 -4 106 96
use mux4_dp_1x  mux4_dp_1x_2
timestamp 1484419186
transform 1 0 0 0 1 550
box -6 -4 106 96
use mux4_dp_1x  mux4_dp_1x_3
timestamp 1484419186
transform 1 0 0 0 1 440
box -6 -4 106 96
use mux4_dp_1x  mux4_dp_1x_4
timestamp 1484419186
transform 1 0 0 0 1 330
box -6 -4 106 96
use mux4_dp_1x  mux4_dp_1x_5
timestamp 1484419186
transform 1 0 0 0 1 220
box -6 -4 106 96
use mux4_dp_1x  mux4_dp_1x_6
timestamp 1484419186
transform 1 0 0 0 1 110
box -6 -4 106 96
use mux4_dp_1x  mux4_dp_1x_7
timestamp 1484419186
transform 1 0 0 0 1 0
box -6 -4 106 96
<< labels >>
rlabel metal2 0 918 4 922 1 s0
rlabel metal2 32 918 36 922 1 s1
rlabel metal2 16 34 20 38 1 d0_0_
rlabel metal2 24 34 28 38 1 d1_0_
rlabel metal2 72 33 76 37 1 d3_0_
rlabel metal2 96 37 100 41 1 y_0_
<< end >>
                                                                                                                                                                                                                                                                                                                                                                      mux4_8_10space.mag                                                                                  0000644 �    Asz0000145 00000000237 13050653540 012125  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1487099744
use mux4_dp_1x  mux4_dp_1x_0
array 0 0 112 0 7 110
timestamp 1484419186
transform 1 0 6 0 1 4
box -6 -4 106 96
<< end >>
                                                                                                                                                                                                                                                                                                                                                                 mux4_8.mag                                                                                          0000644 �    Asz0000145 00000000237 13050653313 010607  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1487099595
use mux4_dp_1x  mux4_dp_1x_0
array 0 0 112 0 7 112
timestamp 1484419186
transform 1 0 6 0 1 4
box -6 -4 106 96
<< end >>
                                                                                                                                                                                                                                                                                                                                                                 mux4_dp_1x.mag                                                                                      0000644 �    Asz0000145 00000013276 13045417656 011476  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1484419186
<< nwell >>
rect -6 40 106 96
<< ntransistor >>
rect 11 7 13 13
rect 16 7 18 13
rect 24 7 26 13
rect 29 7 31 13
rect 37 7 39 13
rect 45 7 47 13
rect 53 7 55 13
rect 58 7 60 13
rect 66 7 68 13
rect 71 7 73 13
rect 93 7 95 14
<< ptransistor >>
rect 11 74 13 83
rect 16 74 18 83
rect 24 74 26 83
rect 29 74 31 83
rect 37 74 39 83
rect 45 74 47 83
rect 53 74 55 83
rect 58 74 60 83
rect 66 74 68 83
rect 71 74 73 83
rect 93 73 95 83
<< ndiffusion >>
rect 6 12 11 13
rect 10 8 11 12
rect 6 7 11 8
rect 13 7 16 13
rect 18 12 24 13
rect 18 8 19 12
rect 23 8 24 12
rect 18 7 24 8
rect 26 7 29 13
rect 31 12 37 13
rect 31 8 32 12
rect 36 8 37 12
rect 31 7 37 8
rect 39 12 45 13
rect 39 8 40 12
rect 44 8 45 12
rect 39 7 45 8
rect 47 12 53 13
rect 47 8 48 12
rect 52 8 53 12
rect 47 7 53 8
rect 55 7 58 13
rect 60 12 66 13
rect 60 8 61 12
rect 65 8 66 12
rect 60 7 66 8
rect 68 7 71 13
rect 73 12 78 13
rect 73 8 74 12
rect 73 7 78 8
rect 88 12 93 14
rect 92 8 93 12
rect 88 7 93 8
rect 95 12 100 14
rect 95 8 96 12
rect 95 7 100 8
<< pdiffusion >>
rect 10 74 11 83
rect 13 74 16 83
rect 18 74 19 83
rect 23 74 24 83
rect 26 74 29 83
rect 31 74 32 83
rect 36 74 37 83
rect 39 74 40 83
rect 44 74 45 83
rect 47 74 48 83
rect 52 74 53 83
rect 55 74 58 83
rect 60 74 61 83
rect 65 74 66 83
rect 68 74 71 83
rect 73 74 74 83
rect 88 82 93 83
rect 92 73 93 82
rect 95 82 100 83
rect 95 73 96 82
<< ndcontact >>
rect 6 8 10 12
rect 19 8 23 12
rect 32 8 36 12
rect 40 8 44 12
rect 48 8 52 12
rect 61 8 65 12
rect 74 8 78 12
rect 88 8 92 12
rect 96 8 100 12
<< pdcontact >>
rect 6 74 10 83
rect 19 74 23 83
rect 32 74 36 83
rect 40 74 44 83
rect 48 74 52 83
rect 61 74 65 83
rect 74 74 78 83
rect 88 73 92 82
rect 96 73 100 82
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
rect 40 -2 44 2
rect 48 -2 52 2
rect 56 -2 60 2
rect 64 -2 68 2
rect 72 -2 76 2
rect 80 -2 84 2
rect 88 -2 92 2
rect 96 -2 100 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
rect 32 88 36 92
rect 40 88 44 92
rect 48 88 52 92
rect 56 88 60 92
rect 64 88 68 92
rect 72 88 76 92
rect 80 88 84 92
rect 88 88 92 92
rect 96 88 100 92
<< polysilicon >>
rect 11 83 13 85
rect 16 83 18 85
rect 24 83 26 85
rect 29 83 31 85
rect 37 83 39 85
rect 45 83 47 85
rect 53 83 55 85
rect 58 83 60 85
rect 66 83 68 85
rect 71 83 73 85
rect 93 83 95 85
rect 11 57 13 74
rect 0 22 2 42
rect 8 30 10 56
rect 16 38 18 74
rect 24 52 26 74
rect 0 20 13 22
rect 11 13 13 20
rect 16 13 18 34
rect 22 50 26 52
rect 22 22 24 50
rect 29 46 31 74
rect 37 53 39 74
rect 45 50 47 74
rect 53 60 55 74
rect 58 73 60 74
rect 58 71 62 73
rect 60 53 62 71
rect 66 59 68 74
rect 71 73 73 74
rect 71 71 78 73
rect 66 57 71 59
rect 60 50 61 53
rect 37 45 39 49
rect 45 48 49 50
rect 37 43 44 45
rect 36 29 38 34
rect 42 29 44 43
rect 47 38 49 48
rect 57 42 58 45
rect 47 35 48 38
rect 56 30 58 42
rect 62 35 64 49
rect 36 27 39 29
rect 42 27 47 29
rect 22 20 26 22
rect 24 13 26 20
rect 29 13 31 26
rect 37 13 39 27
rect 45 13 47 27
rect 53 28 58 30
rect 61 33 64 35
rect 53 13 55 28
rect 61 25 63 33
rect 69 29 71 57
rect 76 46 78 71
rect 84 38 86 56
rect 75 33 76 37
rect 81 36 86 38
rect 58 23 63 25
rect 66 27 71 29
rect 58 13 60 23
rect 66 13 68 27
rect 81 16 83 36
rect 71 14 83 16
rect 93 14 95 73
rect 71 13 73 14
rect 11 5 13 7
rect 16 5 18 7
rect 24 5 26 7
rect 29 5 31 7
rect 37 5 39 7
rect 45 5 47 7
rect 53 5 55 7
rect 58 5 60 7
rect 66 5 68 7
rect 71 5 73 7
rect 93 5 95 7
<< polycontact >>
rect 7 56 11 60
rect 0 42 4 46
rect 14 34 18 38
rect 6 26 10 30
rect 36 49 40 53
rect 51 56 55 60
rect 28 42 32 46
rect 61 49 65 53
rect 24 34 28 38
rect 34 34 38 38
rect 28 26 32 30
rect 53 42 57 46
rect 48 34 52 38
rect 83 56 87 60
rect 75 42 79 46
rect 71 33 75 37
rect 89 27 93 31
<< metal1 >>
rect -2 92 102 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 32 92
rect 36 88 40 92
rect 44 88 48 92
rect 52 88 56 92
rect 60 88 64 92
rect 68 88 72 92
rect 76 88 80 92
rect 84 88 88 92
rect 92 88 96 92
rect 100 88 102 92
rect -2 86 102 88
rect 19 83 23 86
rect 61 83 65 86
rect 6 71 10 74
rect 32 71 36 74
rect 48 71 52 74
rect 74 71 78 74
rect 88 82 92 86
rect 96 82 100 83
rect 6 67 36 71
rect 48 67 78 71
rect 11 56 51 60
rect 55 56 80 60
rect 60 49 61 53
rect 4 42 28 46
rect 32 42 53 46
rect 57 42 75 46
rect 96 41 100 73
rect 38 34 48 38
rect 81 30 89 31
rect 10 26 28 30
rect 44 27 89 30
rect 44 26 85 27
rect 6 16 36 20
rect 6 12 10 16
rect 6 7 10 8
rect 19 12 23 13
rect 19 4 23 8
rect 32 12 36 16
rect 48 16 78 20
rect 32 7 36 8
rect 40 7 44 8
rect 48 12 52 16
rect 48 7 52 8
rect 61 12 65 13
rect 61 4 65 8
rect 74 12 78 16
rect 74 7 78 8
rect 88 12 92 14
rect 88 4 92 8
rect 96 12 100 37
rect 96 7 100 8
rect -2 2 102 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 40 2
rect 44 -2 48 2
rect 52 -2 56 2
rect 60 -2 64 2
rect 68 -2 72 2
rect 76 -2 80 2
rect 84 -2 88 2
rect 92 -2 96 2
rect 100 -2 102 2
rect -2 -4 102 -2
<< m2contact >>
rect 40 74 44 75
rect 40 71 44 74
rect 80 56 83 60
rect 83 56 84 60
rect 32 49 36 53
rect 56 49 60 53
rect 0 42 4 46
rect 16 34 18 38
rect 18 34 20 38
rect 24 34 28 38
rect 48 34 52 38
rect 96 37 100 41
rect 72 33 75 37
rect 75 33 76 37
rect 40 26 44 30
rect 40 12 44 14
rect 40 10 44 12
<< metal2 >>
rect 40 30 44 71
rect 40 14 44 26
rect 40 9 44 10
<< labels >>
rlabel metal1 -1 0 -1 0 3 Gnd!
rlabel m2contact 2 44 2 44 1 s0b
rlabel m2contact 18 36 18 36 1 d0
rlabel m2contact 26 36 26 36 1 d1
rlabel m2contact 34 51 34 51 1 s1
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel m2contact 58 51 58 51 1 d2
rlabel m2contact 82 58 82 58 1 s0
rlabel m2contact 98 39 98 39 1 y
rlabel m2contact 74 35 74 35 1 d3
rlabel m2contact 50 36 50 36 1 s1b
<< end >>
                                                                                                                                                                                                                                                                                                                                  nand2_1x.mag                                                                                        0000644 �    Asz0000145 00000003041 13045420314 011066  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1484411139
<< nwell >>
rect -6 40 26 96
<< ntransistor >>
rect 5 7 7 19
rect 10 7 12 19
<< ptransistor >>
rect 5 71 7 83
rect 13 71 15 83
<< ndiffusion >>
rect 0 17 5 19
rect 4 8 5 17
rect 0 7 5 8
rect 7 7 10 19
rect 12 17 17 19
rect 12 8 13 17
rect 12 7 17 8
<< pdiffusion >>
rect 0 81 5 83
rect 4 72 5 81
rect 0 71 5 72
rect 7 81 13 83
rect 7 72 8 81
rect 12 72 13 81
rect 7 71 13 72
rect 15 81 20 83
rect 15 72 16 81
rect 15 71 20 72
<< ndcontact >>
rect 0 8 4 17
rect 13 8 17 17
<< pdcontact >>
rect 0 72 4 81
rect 8 72 12 81
rect 16 72 20 81
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
<< polysilicon >>
rect 5 83 7 85
rect 13 83 15 85
rect 5 19 7 71
rect 13 42 15 71
rect 10 40 15 42
rect 10 19 12 40
rect 5 5 7 7
rect 10 5 12 7
<< polycontact >>
rect 1 35 5 39
rect 15 51 19 55
<< metal1 >>
rect -2 92 22 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 22 92
rect -2 86 22 88
rect 0 81 4 86
rect 0 71 4 72
rect 8 81 12 83
rect 8 47 12 72
rect 16 81 20 86
rect 16 71 20 72
rect 12 43 17 47
rect 0 17 4 19
rect 0 4 4 8
rect 13 17 17 43
rect 13 7 17 8
rect -2 2 22 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 22 2
rect -2 -4 22 -2
<< m2contact >>
rect 16 51 19 55
rect 19 51 20 55
rect 8 43 12 47
rect 0 35 1 39
rect 1 35 4 39
<< labels >>
rlabel m2contact 1 37 1 37 1 A
rlabel m2contact 10 45 10 45 1 Y
rlabel m2contact 18 53 18 53 1 b
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel metal1 -1 0 -1 0 3 Gnd!
<< end >>
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               NAND2X1.mag                                                                                         0000644 �    Asz0000145 00000002643 13055352531 010504  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1488311641
<< nwell >>
rect -8 48 32 105
<< ntransistor >>
rect 7 6 9 26
rect 12 6 14 26
<< ptransistor >>
rect 7 74 9 94
rect 15 74 17 94
<< ndiffusion >>
rect 2 25 7 26
rect 6 6 7 25
rect 9 6 12 26
rect 14 25 19 26
rect 14 6 15 25
<< pdiffusion >>
rect 2 93 7 94
rect 6 74 7 93
rect 9 93 15 94
rect 9 74 10 93
rect 14 74 15 93
rect 17 93 22 94
rect 17 74 18 93
<< ndcontact >>
rect 2 6 6 25
rect 15 6 19 25
<< pdcontact >>
rect 2 74 6 93
rect 10 74 14 93
rect 18 74 22 93
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 7 33 9 74
rect 6 29 9 33
rect 15 61 17 74
rect 15 57 18 61
rect 15 29 17 57
rect 7 26 9 29
rect 12 27 17 29
rect 12 26 14 27
rect 7 4 9 6
rect 12 4 14 6
<< polycontact >>
rect 2 29 6 33
rect 18 57 22 61
<< metal1 >>
rect -2 102 26 103
rect 2 98 14 102
rect 18 98 26 102
rect -2 97 26 98
rect 2 93 6 97
rect 10 93 14 94
rect 18 93 22 97
rect 2 33 6 37
rect 10 26 14 74
rect 18 53 22 57
rect 2 25 6 26
rect 10 25 19 26
rect 10 23 15 25
rect 2 3 6 6
rect -2 2 26 3
rect 2 -2 14 2
rect 18 -2 26 2
rect -2 -3 26 -2
<< labels >>
flabel metal1 4 100 4 100 4 FreeSans 26 0 0 0 vdd
flabel metal1 12 45 12 45 4 FreeSans 26 0 0 0 Y
flabel metal1 4 0 4 0 4 FreeSans 26 0 0 0 gnd
flabel metal1 4 35 4 35 4 FreeSans 26 0 0 0 A
flabel metal1 20 55 20 55 4 FreeSans 26 0 0 0 B
<< end >>
                                                                                             NAND3X1.mag                                                                                         0000644 �    Asz0000145 00000003526 13055352531 010506  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1488311641
<< nwell >>
rect -8 48 40 105
<< ntransistor >>
rect 7 6 9 36
rect 12 6 14 36
rect 17 6 19 36
<< ptransistor >>
rect 7 74 9 94
rect 15 74 17 94
rect 23 74 25 94
<< ndiffusion >>
rect 2 35 7 36
rect 6 6 7 35
rect 9 6 12 36
rect 14 6 17 36
rect 19 35 24 36
rect 19 6 20 35
<< pdiffusion >>
rect 2 93 7 94
rect 6 74 7 93
rect 9 93 15 94
rect 9 74 10 93
rect 14 74 15 93
rect 17 92 23 94
rect 17 78 18 92
rect 22 78 23 92
rect 17 74 23 78
rect 25 93 30 94
rect 25 74 26 93
<< ndcontact >>
rect 2 6 6 35
rect 20 6 24 35
<< pdcontact >>
rect 2 74 6 93
rect 10 74 14 93
rect 18 78 22 92
rect 26 74 30 93
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 23 94 25 96
rect 7 53 9 74
rect 15 73 17 74
rect 6 49 9 53
rect 7 36 9 49
rect 12 71 17 73
rect 12 36 14 71
rect 23 63 25 74
rect 22 59 25 63
rect 23 39 25 59
rect 17 37 25 39
rect 17 36 19 37
rect 7 4 9 6
rect 12 4 14 6
rect 17 4 19 6
<< polycontact >>
rect 2 49 6 53
rect 18 59 22 63
rect 14 43 18 47
<< metal1 >>
rect -2 102 34 103
rect 2 98 14 102
rect 18 98 34 102
rect -2 97 34 98
rect 2 93 6 97
rect 10 93 14 94
rect 18 92 22 97
rect 18 76 22 78
rect 26 93 30 94
rect 11 73 14 74
rect 26 73 29 74
rect 11 70 29 73
rect 18 63 22 67
rect 26 57 29 70
rect 2 53 6 57
rect 26 53 30 57
rect 10 43 14 47
rect 26 37 29 53
rect 21 36 29 37
rect 2 35 6 36
rect 20 35 29 36
rect 24 34 29 35
rect 2 3 6 6
rect -2 2 34 3
rect 2 -2 14 2
rect 18 -2 34 2
rect -2 -3 34 -2
<< labels >>
flabel metal1 12 45 12 45 4 FreeSans 26 0 0 0 B
flabel metal1 4 100 4 100 4 FreeSans 26 0 0 0 vdd
flabel metal1 4 0 4 0 4 FreeSans 26 0 0 0 gnd
flabel metal1 4 55 4 55 4 FreeSans 26 0 0 0 A
flabel metal1 20 65 20 65 4 FreeSans 26 0 0 0 C
flabel metal1 28 55 28 55 4 FreeSans 26 0 0 0 Y
<< end >>
                                                                                                                                                                          nor2_1x.mag                                                                                         0000644 �    Asz0000145 00000003110 13045420314 010741  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1484411102
<< nwell >>
rect -6 40 26 96
<< ntransistor >>
rect 5 7 7 15
rect 13 7 15 15
<< ptransistor >>
rect 5 67 7 83
rect 10 67 12 83
<< ndiffusion >>
rect 0 13 5 15
rect 4 9 5 13
rect 0 7 5 9
rect 7 13 13 15
rect 7 9 8 13
rect 12 9 13 13
rect 7 7 13 9
rect 15 13 20 15
rect 15 9 16 13
rect 15 7 20 9
<< pdiffusion >>
rect 0 82 5 83
rect 4 68 5 82
rect 0 67 5 68
rect 7 67 10 83
rect 12 82 17 83
rect 12 68 13 82
rect 12 67 17 68
<< ndcontact >>
rect 0 9 4 13
rect 8 9 12 13
rect 16 9 20 13
<< pdcontact >>
rect 0 68 4 82
rect 13 68 17 82
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
<< polysilicon >>
rect 5 83 7 85
rect 10 83 12 85
rect 5 47 7 67
rect 1 43 2 47
rect 6 43 7 47
rect 5 15 7 43
rect 10 44 12 67
rect 10 42 15 44
rect 13 15 15 42
rect 5 5 7 7
rect 13 5 15 7
<< polycontact >>
rect 2 43 6 47
rect 15 26 19 30
<< metal1 >>
rect -2 92 22 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 22 92
rect -2 86 22 88
rect 0 82 4 86
rect 0 67 4 68
rect 13 82 17 83
rect 13 37 17 68
rect 12 33 17 37
rect 0 13 4 15
rect 0 4 4 9
rect 8 13 12 33
rect 8 7 12 9
rect 16 13 20 15
rect 16 4 20 9
rect -2 2 22 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 22 2
rect -2 -4 22 -2
<< m2contact >>
rect 0 43 2 47
rect 2 43 4 47
rect 8 33 12 37
rect 16 26 19 30
rect 19 26 20 30
<< labels >>
rlabel m2contact 2 45 2 45 1 a
rlabel m2contact 10 35 10 35 1 y
rlabel m2contact 18 28 18 28 1 b
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel metal1 -1 0 -1 0 3 Gnd!
<< end >>
                                                                                                                                                                                                                                                                                                                                                                                                                                                        NOR2X1.mag                                                                                          0000644 �    Asz0000145 00000002701 13055352531 010415  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1488311641
<< nwell >>
rect -8 48 32 105
<< ntransistor >>
rect 7 6 9 16
rect 15 6 17 16
<< ptransistor >>
rect 7 54 9 94
rect 12 54 14 94
<< ndiffusion >>
rect 2 15 7 16
rect 6 6 7 15
rect 9 15 15 16
rect 9 6 10 15
rect 14 6 15 15
rect 17 15 22 16
rect 17 6 18 15
<< pdiffusion >>
rect 2 93 7 94
rect 6 54 7 93
rect 9 54 12 94
rect 14 93 19 94
rect 14 54 15 93
<< ndcontact >>
rect 2 6 6 15
rect 10 6 14 15
rect 18 6 22 15
<< pdcontact >>
rect 2 54 6 93
rect 15 54 19 93
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 12 94 14 96
rect 7 23 9 54
rect 12 53 14 54
rect 12 51 17 53
rect 6 19 9 23
rect 7 16 9 19
rect 15 47 18 51
rect 15 16 17 47
rect 7 4 9 6
rect 15 4 17 6
<< polycontact >>
rect 2 19 6 23
rect 18 47 22 51
<< metal1 >>
rect -2 102 26 103
rect 2 98 14 102
rect 18 98 26 102
rect -2 97 26 98
rect 2 93 6 97
rect 15 93 19 94
rect 10 54 15 58
rect 11 37 14 54
rect 18 43 22 47
rect 10 33 14 37
rect 2 23 6 27
rect 11 16 14 33
rect 2 15 6 16
rect 10 15 14 16
rect 18 15 22 16
rect 2 3 6 6
rect 18 3 22 6
rect -2 2 26 3
rect 2 -2 14 2
rect 18 -2 26 2
rect -2 -3 26 -2
<< labels >>
flabel metal1 4 100 4 100 4 FreeSans 26 0 0 0 vdd
flabel metal1 20 45 20 45 4 FreeSans 26 0 0 0 B
flabel metal1 4 0 4 0 4 FreeSans 26 0 0 0 gnd
flabel metal1 12 35 12 35 4 FreeSans 26 0 0 0 Y
flabel metal1 4 25 4 25 4 FreeSans 26 0 0 0 A
<< end >>
                                                               OAI21X1.mag                                                                                         0000644 �    Asz0000145 00000003600 13055352531 010447  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1488311641
<< nwell >>
rect -8 48 34 105
<< ntransistor >>
rect 7 6 9 26
rect 15 6 17 26
rect 23 6 25 26
<< ptransistor >>
rect 7 54 9 94
rect 12 54 14 94
rect 20 74 22 94
<< ndiffusion >>
rect 2 25 7 26
rect 6 6 7 25
rect 9 21 15 26
rect 9 7 10 21
rect 14 7 15 21
rect 9 6 15 7
rect 17 25 23 26
rect 17 6 18 25
rect 22 6 23 25
rect 25 25 30 26
rect 25 6 26 25
<< pdiffusion >>
rect 2 93 7 94
rect 6 54 7 93
rect 9 54 12 94
rect 14 93 20 94
rect 14 54 15 93
rect 19 74 20 93
rect 22 93 27 94
rect 22 74 23 93
<< ndcontact >>
rect 2 6 6 25
rect 10 7 14 21
rect 18 6 22 25
rect 26 6 30 25
<< pdcontact >>
rect 2 54 6 93
rect 15 54 19 93
rect 23 74 27 93
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 12 94 14 96
rect 20 94 22 96
rect 20 65 22 74
rect 7 49 9 54
rect 12 53 14 54
rect 12 51 17 53
rect 4 47 9 49
rect 4 33 6 47
rect 15 43 17 51
rect 14 39 17 43
rect 7 26 9 31
rect 15 26 17 39
rect 23 26 25 63
rect 7 4 9 6
rect 15 4 17 6
rect 23 4 25 6
<< polycontact >>
rect 22 63 26 67
rect 10 39 14 43
rect 6 31 10 35
<< metal1 >>
rect -2 102 34 103
rect 2 98 14 102
rect 18 98 34 102
rect -2 97 34 98
rect 2 93 6 97
rect 15 93 19 94
rect 23 93 27 97
rect 23 57 26 63
rect 19 54 20 57
rect 23 54 30 57
rect 10 43 14 47
rect 17 37 20 54
rect 26 53 30 54
rect 2 36 6 37
rect 2 35 10 36
rect 2 33 6 35
rect 17 33 30 37
rect 3 26 21 28
rect 26 26 29 33
rect 2 25 22 26
rect 10 21 14 22
rect 10 3 14 7
rect 26 25 30 26
rect -2 2 34 3
rect 2 -2 14 2
rect 18 -2 34 2
rect -2 -3 34 -2
<< labels >>
flabel metal1 4 0 4 0 4 FreeSans 26 0 0 0 gnd
flabel metal1 4 100 4 100 4 FreeSans 26 0 0 0 vdd
flabel metal1 4 35 4 35 4 FreeSans 26 0 0 0 A
flabel metal1 12 45 12 45 4 FreeSans 26 0 0 0 B
flabel metal1 28 35 28 35 4 FreeSans 26 0 0 0 Y
flabel metal1 28 55 28 55 4 FreeSans 26 0 0 0 C
<< end >>
                                                                                                                                or2_1x_8.mag                                                                                        0000644 �    Asz0000145 00000003674 13045420054 011032  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1484433330
<< metal2 >>
rect 17 817 21 821
rect 0 808 4 812
rect 24 792 28 796
rect 17 707 21 711
rect 0 698 4 702
rect 24 682 28 686
rect 17 597 21 601
rect 0 588 4 592
rect 24 572 28 576
rect 17 487 21 491
rect 0 478 4 482
rect 24 462 28 466
rect 17 377 21 381
rect 0 368 4 372
rect 24 352 28 356
rect 17 267 21 271
rect 0 258 4 262
rect 24 242 28 246
rect 17 157 21 161
rect 0 148 4 152
rect 24 132 28 136
rect 17 47 21 51
rect 0 38 4 42
rect 24 22 28 26
use or2_1x  or2_1x_0
timestamp 1484419682
transform 1 0 0 0 1 770
box -6 -4 34 96
use or2_1x  or2_1x_1
timestamp 1484419682
transform 1 0 0 0 1 660
box -6 -4 34 96
use or2_1x  or2_1x_2
timestamp 1484419682
transform 1 0 0 0 1 550
box -6 -4 34 96
use or2_1x  or2_1x_3
timestamp 1484419682
transform 1 0 0 0 1 440
box -6 -4 34 96
use or2_1x  or2_1x_4
timestamp 1484419682
transform 1 0 0 0 1 330
box -6 -4 34 96
use or2_1x  or2_1x_5
timestamp 1484419682
transform 1 0 0 0 1 220
box -6 -4 34 96
use or2_1x  or2_1x_6
timestamp 1484419682
transform 1 0 0 0 1 110
box -6 -4 34 96
use or2_1x  or2_1x_7
timestamp 1484419682
transform 1 0 0 0 1 0
box -6 -4 34 96
<< labels >>
rlabel metal2 24 22 28 26 1 b_0_
rlabel metal2 17 47 21 51 1 a_0_
rlabel metal2 0 38 4 42 1 y_0_
rlabel metal2 24 132 28 136 1 b_1_
rlabel metal2 0 148 4 152 1 y_1_
rlabel metal2 17 157 21 161 1 a_1_
rlabel metal2 24 242 28 246 1 b_2_
rlabel metal2 0 258 4 262 1 y_2_
rlabel metal2 17 267 21 271 1 a_2_
rlabel metal2 24 352 28 356 1 b_3_
rlabel metal2 0 368 4 372 1 y_3_
rlabel metal2 17 377 21 381 1 a_3_
rlabel metal2 24 462 28 466 1 b_4_
rlabel metal2 0 478 4 482 1 y_4_
rlabel metal2 17 487 21 491 1 a_4_
rlabel metal2 24 572 28 576 1 b_5_
rlabel metal2 0 588 4 592 1 y_5_
rlabel metal2 17 597 21 601 1 a_5_
rlabel metal2 24 682 28 686 1 b_6_
rlabel metal2 0 698 4 702 1 y_6_
rlabel metal2 17 707 21 711 1 a_6_
rlabel metal2 24 792 28 796 1 b_7_
rlabel metal2 0 808 4 812 1 y_7_
rlabel metal2 17 817 21 821 1 a_7_
<< end >>
                                                                    or2_1x.mag                                                                                          0000644 �    Asz0000145 00000004114 13045420054 010571  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1484419682
<< nwell >>
rect -6 40 34 96
<< ntransistor >>
rect 5 7 7 14
rect 13 7 15 13
rect 21 7 23 13
<< ptransistor >>
rect 5 73 7 83
rect 13 71 15 83
rect 18 71 20 83
<< ndiffusion >>
rect 0 12 5 14
rect 4 8 5 12
rect 0 7 5 8
rect 7 13 12 14
rect 7 12 13 13
rect 7 8 8 12
rect 12 8 13 12
rect 7 7 13 8
rect 15 12 21 13
rect 15 8 16 12
rect 20 8 21 12
rect 15 7 21 8
rect 23 12 28 13
rect 23 8 24 12
rect 23 7 28 8
<< pdiffusion >>
rect 0 82 5 83
rect 4 73 5 82
rect 7 82 13 83
rect 7 73 8 82
rect 12 73 13 82
rect 10 71 13 73
rect 15 71 18 83
rect 20 81 25 83
rect 20 72 21 81
rect 20 71 25 72
<< ndcontact >>
rect 0 8 4 12
rect 8 8 12 12
rect 16 8 20 12
rect 24 8 28 12
<< pdcontact >>
rect 0 73 4 82
rect 8 73 12 82
rect 21 72 25 81
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
<< polysilicon >>
rect 5 83 7 85
rect 13 83 15 85
rect 18 83 20 85
rect 5 41 7 73
rect 13 48 15 71
rect 18 57 20 71
rect 18 55 28 57
rect 5 39 11 41
rect 5 14 7 39
rect 19 34 21 50
rect 13 32 21 34
rect 13 13 15 32
rect 26 26 28 55
rect 25 16 28 22
rect 21 14 28 16
rect 21 13 23 14
rect 5 5 7 7
rect 13 5 15 7
rect 21 5 23 7
<< polycontact >>
rect 15 47 19 51
rect 11 38 15 42
rect 24 22 28 26
<< metal1 >>
rect -2 92 30 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 30 92
rect -2 86 30 88
rect 0 82 4 83
rect 8 82 12 86
rect 21 81 25 83
rect 0 42 4 73
rect 21 59 25 72
rect 21 55 28 59
rect 24 42 28 55
rect 15 38 28 42
rect 0 12 4 38
rect 0 7 4 8
rect 8 12 12 14
rect 8 4 12 8
rect 16 12 20 38
rect 16 7 20 8
rect 24 12 28 13
rect 24 4 28 8
rect -2 2 30 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 30 2
rect -2 -4 30 -2
<< m2contact >>
rect 17 47 19 51
rect 19 47 21 51
rect 0 38 4 42
rect 24 22 28 26
<< metal2 >>
rect 16 47 17 51
<< labels >>
rlabel m2contact 19 49 19 49 1 a
rlabel m2contact 26 24 26 24 1 b
rlabel m2contact 2 40 2 40 1 y
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel metal1 -1 0 -1 0 3 Gnd!
<< end >>
                                                                                                                                                                                                                                                                                                                                                                                                                                                    OR2X1.mag                                                                                           0000644 �    Asz0000145 00000003562 13055352531 010305  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1488311641
<< nwell >>
rect -8 48 40 105
<< ntransistor >>
rect 7 6 9 16
rect 15 6 17 16
rect 23 6 25 16
<< ptransistor >>
rect 7 54 9 94
rect 12 54 14 94
rect 20 74 22 94
<< ndiffusion >>
rect 2 15 7 16
rect 6 6 7 15
rect 9 15 15 16
rect 9 6 10 15
rect 14 6 15 15
rect 17 15 23 16
rect 17 6 18 15
rect 22 6 23 15
rect 25 15 30 16
rect 25 6 26 15
<< pdiffusion >>
rect 2 93 7 94
rect 6 54 7 93
rect 9 54 12 94
rect 14 93 20 94
rect 14 54 15 93
rect 19 74 20 93
rect 22 93 27 94
rect 22 74 23 93
<< ndcontact >>
rect 2 6 6 15
rect 10 6 14 15
rect 18 6 22 15
rect 26 6 30 15
<< pdcontact >>
rect 2 54 6 93
rect 15 54 19 93
rect 23 74 27 93
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 12 94 14 96
rect 20 94 22 96
rect 20 73 22 74
rect 20 71 25 73
rect 7 23 9 54
rect 12 43 14 54
rect 12 41 17 43
rect 15 33 17 41
rect 6 19 9 23
rect 7 16 9 19
rect 15 16 17 29
rect 23 16 25 71
rect 7 4 9 6
rect 15 4 17 6
rect 23 4 25 6
<< polycontact >>
rect 19 47 23 51
rect 14 29 18 33
rect 2 19 6 23
<< metal1 >>
rect -2 102 34 103
rect 2 98 14 102
rect 18 98 34 102
rect -2 97 34 98
rect 2 93 6 94
rect 15 93 19 97
rect 23 93 27 94
rect 24 71 30 74
rect 2 51 6 54
rect 2 48 19 51
rect 27 47 30 71
rect 19 39 22 47
rect 26 43 30 47
rect 10 33 14 37
rect 19 36 24 39
rect 11 29 14 33
rect 2 23 6 27
rect 21 24 24 36
rect 11 21 24 24
rect 11 16 14 21
rect 27 16 30 43
rect 2 15 6 16
rect 10 15 14 16
rect 18 15 22 16
rect 26 15 30 16
rect 2 3 6 6
rect 18 3 22 6
rect -2 2 34 3
rect 2 -2 14 2
rect 18 -2 34 2
rect -2 -3 34 -2
<< labels >>
flabel metal1 28 45 28 45 4 FreeSans 26 0 0 0 Y
flabel metal1 12 35 12 35 4 FreeSans 26 0 0 0 B
flabel metal1 4 100 4 100 4 FreeSans 26 0 0 0 vdd
flabel metal1 4 0 4 0 4 FreeSans 26 0 0 0 gnd
flabel metal1 4 25 4 25 4 FreeSans 26 0 0 0 A
<< end >>
                                                                                                                                              XOR2X1.mag                                                                                          0000644 �    Asz0000145 00000006537 13055352531 010442  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1488311641
<< nwell >>
rect -8 48 64 105
<< ntransistor >>
rect 7 6 9 26
rect 16 6 18 26
rect 21 6 23 26
rect 33 6 35 26
rect 38 6 40 26
rect 47 6 49 26
<< ptransistor >>
rect 7 54 9 94
rect 16 54 18 94
rect 21 54 23 94
rect 33 54 35 94
rect 38 54 40 94
rect 47 54 49 94
<< ndiffusion >>
rect 2 25 7 26
rect 6 6 7 25
rect 9 21 16 26
rect 9 7 10 21
rect 14 7 16 21
rect 9 6 16 7
rect 18 6 21 26
rect 23 22 33 26
rect 23 8 26 22
rect 30 8 33 22
rect 23 6 33 8
rect 35 6 38 26
rect 40 21 47 26
rect 40 7 41 21
rect 45 7 47 21
rect 40 6 47 7
rect 49 25 54 26
rect 49 6 50 25
<< pdiffusion >>
rect 2 93 7 94
rect 6 54 7 93
rect 9 92 16 94
rect 9 63 10 92
rect 14 63 16 92
rect 9 54 16 63
rect 18 54 21 94
rect 23 93 33 94
rect 23 54 26 93
rect 30 54 33 93
rect 35 54 38 94
rect 40 92 47 94
rect 40 63 41 92
rect 45 63 47 92
rect 40 54 47 63
rect 49 93 54 94
rect 49 54 50 93
<< ndcontact >>
rect 2 6 6 25
rect 10 7 14 21
rect 26 8 30 22
rect 41 7 45 21
rect 50 6 54 25
<< pdcontact >>
rect 2 54 6 93
rect 10 63 14 92
rect 26 54 30 93
rect 41 63 45 92
rect 50 54 54 93
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
rect 30 -2 34 2
rect 46 -2 50 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
rect 30 98 34 102
rect 46 98 50 102
<< polysilicon >>
rect 7 94 9 96
rect 16 94 18 96
rect 21 94 23 96
rect 33 94 35 96
rect 38 94 40 96
rect 47 94 49 96
rect 7 37 9 54
rect 16 53 18 54
rect 15 51 18 53
rect 15 47 17 51
rect 7 26 9 33
rect 14 29 16 43
rect 21 39 23 54
rect 33 48 35 54
rect 38 53 40 54
rect 47 53 49 54
rect 38 51 49 53
rect 33 46 40 48
rect 38 37 40 46
rect 47 37 49 51
rect 24 35 32 37
rect 14 27 18 29
rect 16 26 18 27
rect 21 27 22 31
rect 30 29 32 35
rect 47 29 49 33
rect 30 27 35 29
rect 21 26 23 27
rect 33 26 35 27
rect 38 27 49 29
rect 38 26 40 27
rect 47 26 49 27
rect 7 4 9 6
rect 16 4 18 6
rect 21 4 23 6
rect 33 4 35 6
rect 38 4 40 6
rect 47 4 49 6
<< polycontact >>
rect 13 43 17 47
rect 6 33 10 37
rect 20 35 24 39
rect 22 27 26 31
rect 36 33 40 37
rect 46 33 50 37
<< metal1 >>
rect -2 102 58 103
rect 2 98 14 102
rect 18 98 30 102
rect 34 98 46 102
rect 50 98 58 102
rect -2 97 58 98
rect 11 94 15 97
rect 2 93 6 94
rect 10 92 15 94
rect 14 63 15 92
rect 10 61 15 63
rect 24 93 32 94
rect 6 54 11 57
rect 24 54 26 93
rect 30 54 32 93
rect 41 92 46 97
rect 45 63 46 92
rect 41 61 46 63
rect 50 93 54 94
rect 46 54 50 57
rect 27 47 30 54
rect 26 43 30 47
rect 2 33 6 37
rect 10 35 20 38
rect 27 37 30 43
rect 10 34 13 35
rect 27 34 32 37
rect 2 26 11 29
rect 2 25 6 26
rect 29 24 32 34
rect 50 33 54 37
rect 36 31 39 33
rect 46 26 54 29
rect 10 21 15 23
rect 14 7 15 21
rect 10 6 15 7
rect 24 22 32 24
rect 50 25 54 26
rect 24 8 26 22
rect 30 8 32 22
rect 24 6 32 8
rect 41 21 46 23
rect 45 7 46 21
rect 11 3 15 6
rect 41 3 46 7
rect -2 2 58 3
rect 2 -2 14 2
rect 18 -2 30 2
rect 34 -2 46 2
rect 50 -2 58 2
rect -2 -3 58 -2
<< m2contact >>
rect 11 54 15 58
rect 42 54 46 58
rect 17 44 21 48
rect 11 26 15 30
rect 18 27 22 31
rect 35 27 39 31
rect 42 26 46 30
<< metal2 >>
rect 11 30 14 54
rect 18 37 21 44
rect 43 37 46 54
rect 18 34 46 37
rect 15 27 18 30
rect 22 27 35 30
rect 43 30 46 34
<< labels >>
flabel metal1 28 45 28 45 4 FreeSans 26 0 0 0 Y
flabel metal1 4 100 4 100 4 FreeSans 26 0 0 0 vdd
flabel metal1 52 35 52 35 4 FreeSans 26 0 0 0 B
flabel metal1 4 35 4 35 4 FreeSans 26 0 0 0 A
flabel metal1 4 0 4 0 4 FreeSans 26 0 0 0 gnd
<< end >>
                                                                                                                                                                 yzdetect_8.mag                                                                                      0000644 �    Asz0000145 00000003240 13045420314 011537  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   magic
tech scmos
timestamp 1484534894
<< metal1 >>
rect 4 648 8 652
rect -4 593 13 597
rect 12 538 16 542
rect -4 373 3 377
rect 17 356 24 360
rect 12 208 16 212
rect 9 153 24 157
rect 4 98 8 102
<< m2contact >>
rect 0 648 4 652
rect 8 648 12 652
rect -8 593 -4 597
rect 8 538 12 542
rect 16 538 20 542
rect -8 373 -4 377
rect 24 356 28 360
rect 8 208 12 212
rect 16 208 20 212
rect 24 153 28 157
rect 0 98 4 102
rect 8 98 12 102
<< metal2 >>
rect 0 703 4 707
rect 8 652 12 696
rect 16 686 20 690
rect -8 377 -4 593
rect 0 586 4 648
rect 16 542 20 604
rect 0 483 4 487
rect 8 474 12 538
rect 16 466 20 470
rect 8 363 12 367
rect 0 263 4 267
rect 8 212 12 256
rect 16 246 20 250
rect 16 162 20 208
rect 24 157 28 356
rect 0 102 4 145
rect 0 43 4 47
rect 8 34 12 98
rect 16 26 20 30
use nor2_1x  nor2_1x_0
timestamp 1484411102
transform 1 0 0 0 1 660
box -6 -4 26 96
use nand2_1x  nand2_1x_0
timestamp 1484411139
transform 1 0 0 0 1 550
box -6 -4 26 96
use nor2_1x  nor2_1x_1
timestamp 1484411102
transform 1 0 0 0 1 440
box -6 -4 26 96
use nor2_1x  nor2_1x_2
timestamp 1484411102
transform 1 0 0 0 1 330
box -6 -4 26 96
use nor2_1x  nor2_1x_3
timestamp 1484411102
transform 1 0 0 0 1 220
box -6 -4 26 96
use nand2_1x  nand2_1x_1
timestamp 1484411139
transform 1 0 0 0 1 110
box -6 -4 26 96
use nor2_1x  nor2_1x_4
timestamp 1484411102
transform 1 0 0 0 1 0
box -6 -4 26 96
<< labels >>
rlabel metal2 16 26 20 30 1 a_1_
rlabel metal2 0 43 4 47 1 a_0_
rlabel metal2 0 263 4 267 1 a_2_
rlabel metal2 16 246 20 250 1 a_3_
rlabel metal2 8 363 12 367 1 zero
rlabel metal2 0 483 4 487 1 a_4_
rlabel metal2 16 466 20 470 1 a_5_
rlabel metal2 16 686 20 690 1 a_7_
rlabel metal2 0 703 4 707 1 a_6_
<< end >>
                                                                                                                                                                                                                                                                                                                                                                basic-test.irsim                                                                                    0000644 �    Asz0000145 00000007721 13055367521 012115  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   ﻿# Basic IRSIM test file shell for ECE 425 Lab 4.

# In order to ensure that your layout will be testable by the instructors,
# make sure that you can source this file without any errors, especially
# errors for unknown node names.  The remainder of the file may or may not
# be useful for your own testing.


# Basic setup.
l Gnd!
h Vdd!
l less
stepsize 100
logfile alu.log

# Set up the vectors.
vector funct funct_5 funct_4 funct_3 funct_2 funct_1 funct_0
vector alu_op alu_op_1 alu_op_0
vector op op6 op5 op4 op3 op2 op1 op0
vector a a7 a6 a5 a4 a3 a2 a1 a0
vector b b7 b6 b5 b4 b3 b2 b1 b0
vector result result7 result6 result5 result4 result3 result2 result1 result0

# Add the top-level signals to the watch list.  This causes theie values to be
# displayed after each step.
w funct alu_op a b result op


#
# A sample test; you will need a few more ...
#

# AND1
setvector funct 100100
setvector alu_op 10
setvector a 01010101
setvector b 11111111
s
assert result 01010101

# AND2
setvector funct 100100
setvector alu_op 10
setvector a 01010101
setvector b 10101010
s
assert result 00000000

# AND3
setvector funct 100100
setvector alu_op 10
setvector a 11111001
setvector b 00001001
s
assert result 00001001


# OR1
setvector funct 100101
setvector alu_op 10
setvector a 01010101
setvector b 11111111
s
assert result 11111111

# OR2
setvector funct 100101
setvector alu_op 10
setvector a 01010101
setvector b 00000010
s
assert result 01010111

# OR3
setvector funct 100101
setvector alu_op 10
setvector a 00001111
setvector b 11001111
s
assert result 11001111

# NOR1
setvector funct 100111
setvector alu_op 10
setvector a 00001111
setvector b 11001111
s
assert result 00110000

# NOR2
setvector funct 100111
setvector alu_op 10
setvector a 01010101
setvector b 00000010
s
assert result 10101000

# NOR3
setvector funct 100111
setvector alu_op 10
setvector a 00001111
setvector b 11111111
s
assert result 00000000

# XOR1
setvector funct 100110
setvector alu_op 10
setvector a 01010101
setvector b 11111111
s
assert result 10101010

# XOR2
setvector funct 100110
setvector alu_op 10
setvector a 01010101
setvector b 11110000
s
assert result 10100101

# XOR3
setvector funct 100110
setvector alu_op 10
setvector a 11110000
setvector b 11111111
s
assert result 00001111

# ADD1
setvector funct 100000
setvector alu_op 10
setvector a 01110000
setvector b 01111111
s
assert result 11101111

# ADD2
setvector funct 100000
setvector alu_op 10
setvector a 00001010
setvector b 01101000
s
assert result 01110010

# ADD3
setvector funct 100000
setvector alu_op 10
setvector a 00001010
setvector b 01111111
s
assert result 10001001

# sub1
setvector funct 100010
setvector alu_op 10
setvector a 01111111
setvector b 00001010
s
assert result 01110101

# sub2
setvector funct 100010
setvector alu_op 10
setvector a 00001111
setvector b 00001010
s
assert result 00000101

# sub3
setvector funct 100010
setvector alu_op 10
setvector a 01111000
setvector b 00001010
s
assert result 01101110

# SLT1
setvector funct 101011
setvector alu_op 10
setvector a 01111000
setvector b 00001010
s
assert result 00000000

# SLT2
setvector funct 101011
setvector alu_op 10
setvector a 00001111
setvector b 00001010
s
assert result 00000000

# SLT3
setvector funct 101011
setvector alu_op 10
setvector a 00000000
setvector b 00001010
s
assert result 00000001

# SLT4
setvector funct 101011
setvector alu_op 10
setvector a 00000101
setvector b 00101010
s
assert result 00000001

# SLT5
setvector funct 101011
setvector alu_op 10
setvector a 11111111
setvector b 00000000
s
assert result 00000000

# SLT6
setvector funct 101011
setvector alu_op 10
setvector a 00000000
setvector b 11111111
s
assert result 00000001

# SLT7
setvector funct 101011
setvector alu_op 10
setvector a 11111110
setvector b 11111111
s
assert result 00000001

# SLT8
setvector funct 101011
setvector alu_op 10
setvector a 11111111
setvector b 11111111
s
assert result 00000000

# SLT9
setvector funct 101011
setvector alu_op 10
setvector a 00000000
setvector b 00000000
s
assert result 00000000
                                               alt_alu_with_ctl.sim                                                                                0000644 �    Asz0000145 00000233550 13055370467 013046  0                                                                                                    ustar   hany                                                                                                                                                                                                                                                   | units: 30 tech: scmos format: MIT
p alu_ctl_0/NOR2X1_0/B Vdd! alu_ctl_0/NOR2X1_2/a_9_54# 2 40 673 144
p funct_3 alu_ctl_0/NOR2X1_2/a_9_54# alu_ctl_0/NOR2X1_2/Y 2 40 678 144
n alu_ctl_0/NOR2X1_0/B Gnd! alu_ctl_0/NOR2X1_2/Y 2 10 673 96
n funct_3 alu_ctl_0/NOR2X1_2/Y Gnd! 2 10 681 96
p alu_ctl_0/NOR2X1_1/Y Vdd! alu_ctl_0/NOR2X1_0/B 2 20 649 164
p funct_5 alu_ctl_0/NOR2X1_0/B Vdd! 2 20 657 164
n alu_ctl_0/NOR2X1_1/Y Gnd! alu_ctl_0/NAND2X1_6/a_9_6# 2 20 649 96
n funct_5 alu_ctl_0/NAND2X1_6/a_9_6# alu_ctl_0/NOR2X1_0/B 2 20 654 96
p funct_4 Vdd! alu_ctl_0/NOR2X1_1/a_9_54# 2 40 593 144
p alu_op_0 alu_ctl_0/NOR2X1_1/a_9_54# alu_ctl_0/NOR2X1_1/Y 2 40 598 144
n funct_4 Gnd! alu_ctl_0/NOR2X1_1/Y 2 10 593 96
n alu_op_0 alu_ctl_0/NOR2X1_1/Y Gnd! 2 10 601 96
p alu_ctl_0/NOR2X1_0/A Vdd! alu_ctl_0/NOR2X1_0/a_9_54# 2 40 561 144
p alu_ctl_0/NOR2X1_0/B alu_ctl_0/NOR2X1_0/a_9_54# alu_ctl_0/NOR2X1_0/Y 2 40 566 144
n alu_ctl_0/NOR2X1_0/A Gnd! alu_ctl_0/NOR2X1_0/Y 2 10 561 96
n alu_ctl_0/NOR2X1_0/B alu_ctl_0/NOR2X1_0/Y Gnd! 2 10 569 96
p alu_ctl_0/OAI21X1_7/A Vdd! alu_ctl_0/OAI21X1_7/a_9_54# 2 40 506 144
p alu_ctl_0/OAI21X1_7/B alu_ctl_0/OAI21X1_7/a_9_54# op6 2 40 501 144
p alu_ctl_0/INVX2_0/Y op6 Vdd! 2 20 493 164
n alu_ctl_0/OAI21X1_7/A alu_ctl_0/OAI21X1_7/a_2_6# Gnd! 2 20 506 96
n alu_ctl_0/OAI21X1_7/B Gnd! alu_ctl_0/OAI21X1_7/a_2_6# 2 20 498 96
n alu_ctl_0/INVX2_0/Y alu_ctl_0/OAI21X1_7/a_2_6# op6 2 20 490 96
p alu_ctl_0/NOR2X1_2/Y Vdd! alu_ctl_0/OAI21X1_6/C 2 20 657 215
p alu_ctl_0/NAND2X1_5/B alu_ctl_0/OAI21X1_6/C Vdd! 2 20 665 215
n alu_ctl_0/NOR2X1_2/Y Gnd! alu_ctl_0/NAND2X1_5/a_9_6# 2 20 657 283
n alu_ctl_0/NAND2X1_5/B alu_ctl_0/NAND2X1_5/a_9_6# alu_ctl_0/OAI21X1_6/C 2 20 662 283
p alu_op_1 Vdd! alu_ctl_0/OAI21X1_6/a_9_54# 2 40 609 235
p alu_op_0 alu_ctl_0/OAI21X1_6/a_9_54# op5 2 40 614 235
p alu_ctl_0/OAI21X1_6/C op5 Vdd! 2 20 622 215
n alu_op_1 alu_ctl_0/OAI21X1_6/a_2_6# Gnd! 2 20 609 283
n alu_op_0 Gnd! alu_ctl_0/OAI21X1_6/a_2_6# 2 20 617 283
n alu_ctl_0/OAI21X1_6/C alu_ctl_0/OAI21X1_6/a_2_6# op5 2 20 625 283
p alu_ctl_0/NOR2X1_2/Y Vdd! alu_ctl_0/INVX2_3/A 2 20 594 215
p alu_op_1 alu_ctl_0/INVX2_3/A Vdd! 2 20 586 215
n alu_ctl_0/NOR2X1_2/Y Gnd! alu_ctl_0/NAND2X1_4/a_9_6# 2 20 594 283
n alu_op_1 alu_ctl_0/NAND2X1_4/a_9_6# alu_ctl_0/INVX2_3/A 2 20 589 283
p alu_ctl_0/NOR2X1_0/A Vdd! alu_ctl_0/NAND3X1_2/Y 2 20 554 215
p alu_ctl_0/INVX2_5/Y alu_ctl_0/NAND3X1_2/Y Vdd! 2 20 546 215
p alu_ctl_0/NOR2X1_2/Y Vdd! alu_ctl_0/NAND3X1_2/Y 2 20 538 215
n alu_ctl_0/NOR2X1_0/A Gnd! alu_ctl_0/NAND3X1_2/a_9_6# 2 30 554 283
n alu_ctl_0/INVX2_5/Y alu_ctl_0/NAND3X1_2/a_9_6# alu_ctl_0/NAND3X1_2/a_14_6# 2 30 549 283
n alu_ctl_0/NOR2X1_2/Y alu_ctl_0/NAND3X1_2/a_14_6# alu_ctl_0/NAND3X1_2/Y 2 30 544 283
p funct_0 Vdd! alu_ctl_0/NOR2X1_0/A 2 20 481 215
p alu_ctl_0/INVX2_2/Y alu_ctl_0/NOR2X1_0/A Vdd! 2 20 489 215
n funct_0 Gnd! alu_ctl_0/NAND2X1_3/a_9_6# 2 20 481 283
n alu_ctl_0/INVX2_2/Y alu_ctl_0/NAND2X1_3/a_9_6# alu_ctl_0/NOR2X1_0/A 2 20 486 283
p alu_ctl_0/INVX2_6/A Vdd! alu_ctl_0/INVX2_6/Y 2 40 689 344
n alu_ctl_0/INVX2_6/A Gnd! alu_ctl_0/INVX2_6/Y 2 20 689 296
p alu_ctl_0/INVX2_5/Y Vdd! alu_ctl_0/OAI21X1_5/a_9_54# 2 40 617 344
p funct_0 alu_ctl_0/OAI21X1_5/a_9_54# alu_ctl_0/INVX2_6/A 2 40 622 344
p alu_ctl_0/NAND3X1_0/Y alu_ctl_0/INVX2_6/A Vdd! 2 20 630 364
n alu_ctl_0/INVX2_5/Y alu_ctl_0/OAI21X1_5/a_2_6# Gnd! 2 20 617 296
n funct_0 Gnd! alu_ctl_0/OAI21X1_5/a_2_6# 2 20 625 296
n alu_ctl_0/NAND3X1_0/Y alu_ctl_0/OAI21X1_5/a_2_6# alu_ctl_0/INVX2_6/A 2 20 633 296
p alu_ctl_0/NOR2X1_0/Y Vdd! alu_ctl_0/INVX2_1/A 2 20 562 364
p alu_op_1 alu_ctl_0/INVX2_1/A Vdd! 2 20 554 364
p alu_ctl_0/AND2X2_0/Y Vdd! alu_ctl_0/INVX2_1/A 2 20 546 364
n alu_ctl_0/NOR2X1_0/Y Gnd! alu_ctl_0/NAND3X1_1/a_9_6# 2 30 562 296
n alu_op_1 alu_ctl_0/NAND3X1_1/a_9_6# alu_ctl_0/NAND3X1_1/a_14_6# 2 30 557 296
n alu_ctl_0/AND2X2_0/Y alu_ctl_0/NAND3X1_1/a_14_6# alu_ctl_0/INVX2_1/A 2 30 552 296
p funct_1 Vdd! alu_ctl_0/OAI21X1_7/A 2 20 489 364
p funct_0 alu_ctl_0/OAI21X1_7/A Vdd! 2 20 497 364
n funct_1 Gnd! alu_ctl_0/NAND2X1_2/a_9_6# 2 20 489 296
n funct_0 alu_ctl_0/NAND2X1_2/a_9_6# alu_ctl_0/OAI21X1_7/A 2 20 494 296
p funct_1 Vdd! alu_ctl_0/INVX2_5/Y 2 40 473 344
n funct_1 Gnd! alu_ctl_0/INVX2_5/Y 2 20 473 296
p funct_0 Vdd! alu_ctl_0/OAI21X1_4/a_9_54# 2 40 657 435
p alu_ctl_0/XOR2X1_0/Y alu_ctl_0/OAI21X1_4/a_9_54# alu_ctl_0/NAND2X1_5/B 2 40 662 435
p alu_ctl_0/NAND3X1_0/Y alu_ctl_0/NAND2X1_5/B Vdd! 2 20 670 415
n funct_0 alu_ctl_0/OAI21X1_4/a_2_6# Gnd! 2 20 657 483
n alu_ctl_0/XOR2X1_0/Y Gnd! alu_ctl_0/OAI21X1_4/a_2_6# 2 20 665 483
n alu_ctl_0/NAND3X1_0/Y alu_ctl_0/OAI21X1_4/a_2_6# alu_ctl_0/NAND2X1_5/B 2 20 673 483
p funct_0 Vdd! alu_ctl_0/NAND3X1_0/Y 2 20 593 415
p alu_ctl_0/INVX2_5/Y alu_ctl_0/NAND3X1_0/Y Vdd! 2 20 601 415
p funct_2 Vdd! alu_ctl_0/NAND3X1_0/Y 2 20 609 415
n funct_0 Gnd! alu_ctl_0/NAND3X1_0/a_9_6# 2 30 593 483
n alu_ctl_0/INVX2_5/Y alu_ctl_0/NAND3X1_0/a_9_6# alu_ctl_0/NAND3X1_0/a_14_6# 2 30 598 483
n funct_2 alu_ctl_0/NAND3X1_0/a_14_6# alu_ctl_0/NAND3X1_0/Y 2 30 603 483
p alu_op_1 Vdd! alu_ctl_0/INVX2_4/Y 2 40 482 435
n alu_op_1 Gnd! alu_ctl_0/INVX2_4/Y 2 20 482 483
p funct_1 Vdd! alu_ctl_0/AND2X2_0/a_2_6# 2 20 674 564
p funct_3 alu_ctl_0/AND2X2_0/a_2_6# Vdd! 2 20 666 564
p alu_ctl_0/AND2X2_0/a_2_6# Vdd! alu_ctl_0/AND2X2_0/Y 2 40 658 544
n funct_1 alu_ctl_0/AND2X2_0/a_2_6# alu_ctl_0/AND2X2_0/a_9_6# 2 20 674 496
n funct_3 alu_ctl_0/AND2X2_0/a_9_6# Gnd! 2 20 669 496
n alu_ctl_0/AND2X2_0/a_2_6# Gnd! alu_ctl_0/AND2X2_0/Y 2 20 661 496
p funct_2 Vdd! alu_ctl_0/OAI21X1_7/B 2 20 586 564
p alu_ctl_0/INVX2_3/Y alu_ctl_0/OAI21X1_7/B Vdd! 2 20 578 564
n funct_2 Gnd! alu_ctl_0/NAND2X1_1/a_9_6# 2 20 586 496
n alu_ctl_0/INVX2_3/Y alu_ctl_0/NAND2X1_1/a_9_6# alu_ctl_0/OAI21X1_7/B 2 20 581 496
p funct_0 alu_ctl_0/OR2X1_0/a_2_54# alu_ctl_0/OR2X1_0/a_9_54# 2 40 514 544
p funct_2 alu_ctl_0/OR2X1_0/a_9_54# Vdd! 2 40 509 544
p alu_ctl_0/OR2X1_0/a_2_54# Vdd! alu_ctl_0/OR2X1_0/Y 2 20 501 564
n funct_0 Gnd! alu_ctl_0/OR2X1_0/a_2_54# 2 10 514 496
n funct_2 alu_ctl_0/OR2X1_0/a_2_54# Gnd! 2 10 506 496
n alu_ctl_0/OR2X1_0/a_2_54# Gnd! alu_ctl_0/OR2X1_0/Y 2 10 498 496
p alu_ctl_0/INVX2_6/Y Vdd! alu_ctl_0/OAI21X1_3/a_9_54# 2 40 666 635
p alu_ctl_0/INVX2_3/A alu_ctl_0/OAI21X1_3/a_9_54# op4 2 40 661 635
p alu_ctl_0/OAI21X1_2/C op4 Vdd! 2 20 653 615
n alu_ctl_0/INVX2_6/Y alu_ctl_0/OAI21X1_3/a_2_6# Gnd! 2 20 666 683
n alu_ctl_0/INVX2_3/A Gnd! alu_ctl_0/OAI21X1_3/a_2_6# 2 20 658 683
n alu_ctl_0/OAI21X1_2/C alu_ctl_0/OAI21X1_3/a_2_6# op4 2 20 650 683
p alu_ctl_0/INVX2_3/Y Vdd! alu_ctl_0/OAI21X1_2/B 2 20 594 615
p funct_1 alu_ctl_0/OAI21X1_2/B Vdd! 2 20 586 615
n alu_ctl_0/INVX2_3/Y Gnd! alu_ctl_0/NAND2X1_0/a_9_6# 2 20 594 683
n funct_1 alu_ctl_0/NAND2X1_0/a_9_6# alu_ctl_0/OAI21X1_2/B 2 20 589 683
p alu_ctl_0/INVX2_3/A Vdd! alu_ctl_0/INVX2_3/Y 2 40 570 635
n alu_ctl_0/INVX2_3/A Gnd! alu_ctl_0/INVX2_3/Y 2 20 570 683
p alu_ctl_0/OR2X1_0/Y Vdd! alu_ctl_0/OAI21X1_2/a_9_54# 2 40 506 635
p alu_ctl_0/OAI21X1_2/B alu_ctl_0/OAI21X1_2/a_9_54# op2 2 40 501 635
p alu_ctl_0/OAI21X1_2/C op2 Vdd! 2 20 493 615
n alu_ctl_0/OR2X1_0/Y alu_ctl_0/OAI21X1_2/a_2_6# Gnd! 2 20 506 683
n alu_ctl_0/OAI21X1_2/B Gnd! alu_ctl_0/OAI21X1_2/a_2_6# 2 20 498 683
n alu_ctl_0/OAI21X1_2/C alu_ctl_0/OAI21X1_2/a_2_6# op2 2 20 490 683
p funct_2 Vdd! alu_ctl_0/INVX2_2/Y 2 40 690 744
n funct_2 Gnd! alu_ctl_0/INVX2_2/Y 2 20 690 696
p funct_2 alu_ctl_0/XOR2X1_0/a_2_6# Vdd! 2 40 633 744
p alu_ctl_0/XOR2X1_0/a_13_43# Vdd! alu_ctl_0/XOR2X1_0/a_18_54# 2 40 642 744
p funct_2 alu_ctl_0/XOR2X1_0/a_18_54# alu_ctl_0/XOR2X1_0/Y 2 40 647 744
p alu_ctl_0/XOR2X1_0/a_2_6# alu_ctl_0/XOR2X1_0/Y alu_ctl_0/XOR2X1_0/a_35_54# 2 40 659 744
p funct_1 alu_ctl_0/XOR2X1_0/a_35_54# Vdd! 2 40 664 744
p funct_1 Vdd! alu_ctl_0/XOR2X1_0/a_13_43# 2 40 673 744
n funct_2 alu_ctl_0/XOR2X1_0/a_2_6# Gnd! 2 20 633 696
n alu_ctl_0/XOR2X1_0/a_13_43# Gnd! alu_ctl_0/XOR2X1_0/a_18_6# 2 20 642 696
n alu_ctl_0/XOR2X1_0/a_2_6# alu_ctl_0/XOR2X1_0/a_18_6# alu_ctl_0/XOR2X1_0/Y 2 20 647 696
n funct_2 alu_ctl_0/XOR2X1_0/Y alu_ctl_0/XOR2X1_0/a_35_6# 2 20 659 696
n funct_1 alu_ctl_0/XOR2X1_0/a_35_6# Gnd! 2 20 664 696
n funct_1 Gnd! alu_ctl_0/XOR2X1_0/a_13_43# 2 20 673 696
p alu_ctl_0/INVX2_3/A Vdd! alu_ctl_0/OAI21X1_1/a_9_54# 2 40 585 744
p alu_ctl_0/INVX2_2/Y alu_ctl_0/OAI21X1_1/a_9_54# op0 2 40 590 744
p alu_ctl_0/INVX2_1/A op0 Vdd! 2 20 598 764
n alu_ctl_0/INVX2_3/A alu_ctl_0/OAI21X1_1/a_2_6# Gnd! 2 20 585 696
n alu_ctl_0/INVX2_2/Y Gnd! alu_ctl_0/OAI21X1_1/a_2_6# 2 20 593 696
n alu_ctl_0/INVX2_1/A alu_ctl_0/OAI21X1_1/a_2_6# op0 2 20 601 696
p alu_op_1 Vdd! alu_ctl_0/OAI21X1_0/a_9_54# 2 40 505 744
p alu_op_0 alu_ctl_0/OAI21X1_0/a_9_54# op3 2 40 510 744
p alu_ctl_0/NAND3X1_2/Y op3 Vdd! 2 20 518 764
n alu_op_1 alu_ctl_0/OAI21X1_0/a_2_6# Gnd! 2 20 505 696
n alu_op_0 Gnd! alu_ctl_0/OAI21X1_0/a_2_6# 2 20 513 696
n alu_ctl_0/NAND3X1_2/Y alu_ctl_0/OAI21X1_0/a_2_6# op3 2 20 521 696
p alu_ctl_0/INVX2_1/A Vdd! op1 2 40 650 835
n alu_ctl_0/INVX2_1/A Gnd! op1 2 20 650 883
p alu_ctl_0/INVX2_4/Y alu_ctl_0/AOI21X1_0/a_2_54# Vdd! 2 40 553 835
p alu_op_0 Vdd! alu_ctl_0/AOI21X1_0/a_2_54# 2 40 561 835
p op1 alu_ctl_0/AOI21X1_0/a_2_54# alu_ctl_0/OAI21X1_2/C 2 40 569 835
n alu_ctl_0/INVX2_4/Y Gnd! alu_ctl_0/AOI21X1_0/a_12_6# 2 20 556 883
n alu_op_0 alu_ctl_0/AOI21X1_0/a_12_6# alu_ctl_0/OAI21X1_2/C 2 20 561 883
n op1 alu_ctl_0/OAI21X1_2/C Gnd! 2 10 569 883
p op2 Vdd! alu_ctl_0/INVX2_0/Y 2 40 481 835
n op2 Gnd! alu_ctl_0/INVX2_0/Y 2 20 481 883
p mux3_1x_8_0/mux3_dp_1x_7/s0 mux3_1x_8_0/mux3_dp_1x_7/a_0_74# mux3_1x_8_0/mux3_dp_1x_7/a_7_74# 2 9 301 78
p adder_8_0/s_0_ mux3_1x_8_0/mux3_dp_1x_7/a_7_74# Vdd! 2 9 306 78
p muxy7 Vdd! mux3_1x_8_0/mux3_dp_1x_7/a_20_74# 2 9 314 78
p mux3_1x_8_0/mux3_dp_1x_7/s0b mux3_1x_8_0/mux3_dp_1x_7/a_20_74# mux3_1x_8_0/mux3_dp_1x_7/a_0_74# 2 9 319 78
p mux3_1x_8_0/mux3_dp_1x_7/s1 mux3_1x_8_0/mux3_dp_1x_7/a_0_74# mux3_1x_8_0/mux3_dp_1x_7/a_33_7# 2 9 327 78
p mux3_1x_8_0/mux3_dp_1x_7/s1b mux3_1x_8_0/mux3_dp_1x_7/a_33_7# mux3_1x_8_0/mux3_dp_1x_7/a_41_74# 2 9 335 78
p inv_1x_0/y mux3_1x_8_0/mux3_dp_1x_7/a_41_74# Vdd! 2 9 340 78
p mux3_1x_8_0/mux3_dp_1x_7/a_33_7# result0 Vdd! 2 10 355 77
n mux3_1x_8_0/mux3_dp_1x_7/s0 mux3_1x_8_0/mux3_dp_1x_7/a_0_7# mux3_1x_8_0/mux3_dp_1x_7/a_7_7# 2 6 301 11
n muxy7 mux3_1x_8_0/mux3_dp_1x_7/a_7_7# Gnd! 2 6 306 11
n adder_8_0/s_0_ Gnd! mux3_1x_8_0/mux3_dp_1x_7/a_20_7# 2 6 314 11
n mux3_1x_8_0/mux3_dp_1x_7/s0b mux3_1x_8_0/mux3_dp_1x_7/a_20_7# mux3_1x_8_0/mux3_dp_1x_7/a_0_7# 2 6 319 11
n mux3_1x_8_0/mux3_dp_1x_7/s1b mux3_1x_8_0/mux3_dp_1x_7/a_0_7# mux3_1x_8_0/mux3_dp_1x_7/a_33_7# 2 6 327 11
n mux3_1x_8_0/mux3_dp_1x_7/s1 mux3_1x_8_0/mux3_dp_1x_7/a_33_7# mux3_1x_8_0/mux3_dp_1x_7/a_41_7# 2 6 335 11
n inv_1x_0/y mux3_1x_8_0/mux3_dp_1x_7/a_41_7# Gnd! 2 6 340 11
n mux3_1x_8_0/mux3_dp_1x_7/a_33_7# Gnd! result0 2 7 358 16
p mux3_1x_8_0/mux3_dp_1x_7/s0 mux3_1x_8_0/mux3_dp_1x_6/a_0_74# mux3_1x_8_0/mux3_dp_1x_6/a_7_74# 2 9 301 188
p adder_8_0/s_1_ mux3_1x_8_0/mux3_dp_1x_6/a_7_74# Vdd! 2 9 306 188
p adder_8_0/b_1_ Vdd! mux3_1x_8_0/mux3_dp_1x_6/a_20_74# 2 9 314 188
p mux3_1x_8_0/mux3_dp_1x_7/s0b mux3_1x_8_0/mux3_dp_1x_6/a_20_74# mux3_1x_8_0/mux3_dp_1x_6/a_0_74# 2 9 319 188
p mux3_1x_8_0/mux3_dp_1x_7/s1 mux3_1x_8_0/mux3_dp_1x_6/a_0_74# mux3_1x_8_0/mux3_dp_1x_6/a_33_7# 2 9 327 188
p mux3_1x_8_0/mux3_dp_1x_7/s1b mux3_1x_8_0/mux3_dp_1x_6/a_33_7# mux3_1x_8_0/mux3_dp_1x_6/a_41_74# 2 9 335 188
p less mux3_1x_8_0/mux3_dp_1x_6/a_41_74# Vdd! 2 9 340 188
p mux3_1x_8_0/mux3_dp_1x_6/a_33_7# result1 Vdd! 2 10 355 187
n mux3_1x_8_0/mux3_dp_1x_7/s0 mux3_1x_8_0/mux3_dp_1x_6/a_0_7# mux3_1x_8_0/mux3_dp_1x_6/a_7_7# 2 6 301 121
n adder_8_0/b_1_ mux3_1x_8_0/mux3_dp_1x_6/a_7_7# Gnd! 2 6 306 121
n adder_8_0/s_1_ Gnd! mux3_1x_8_0/mux3_dp_1x_6/a_20_7# 2 6 314 121
n mux3_1x_8_0/mux3_dp_1x_7/s0b mux3_1x_8_0/mux3_dp_1x_6/a_20_7# mux3_1x_8_0/mux3_dp_1x_6/a_0_7# 2 6 319 121
n mux3_1x_8_0/mux3_dp_1x_7/s1b mux3_1x_8_0/mux3_dp_1x_6/a_0_7# mux3_1x_8_0/mux3_dp_1x_6/a_33_7# 2 6 327 121
n mux3_1x_8_0/mux3_dp_1x_7/s1 mux3_1x_8_0/mux3_dp_1x_6/a_33_7# mux3_1x_8_0/mux3_dp_1x_6/a_41_7# 2 6 335 121
n less mux3_1x_8_0/mux3_dp_1x_6/a_41_7# Gnd! 2 6 340 121
n mux3_1x_8_0/mux3_dp_1x_6/a_33_7# Gnd! result1 2 7 358 126
p mux3_1x_8_0/mux3_dp_1x_7/s0 mux3_1x_8_0/mux3_dp_1x_5/a_0_74# mux3_1x_8_0/mux3_dp_1x_5/a_7_74# 2 9 301 298
p adder_8_0/s_2_ mux3_1x_8_0/mux3_dp_1x_5/a_7_74# Vdd! 2 9 306 298
p adder_8_0/b_2_ Vdd! mux3_1x_8_0/mux3_dp_1x_5/a_20_74# 2 9 314 298
p mux3_1x_8_0/mux3_dp_1x_7/s0b mux3_1x_8_0/mux3_dp_1x_5/a_20_74# mux3_1x_8_0/mux3_dp_1x_5/a_0_74# 2 9 319 298
p mux3_1x_8_0/mux3_dp_1x_7/s1 mux3_1x_8_0/mux3_dp_1x_5/a_0_74# mux3_1x_8_0/mux3_dp_1x_5/a_33_7# 2 9 327 298
p mux3_1x_8_0/mux3_dp_1x_7/s1b mux3_1x_8_0/mux3_dp_1x_5/a_33_7# mux3_1x_8_0/mux3_dp_1x_5/a_41_74# 2 9 335 298
p less mux3_1x_8_0/mux3_dp_1x_5/a_41_74# Vdd! 2 9 340 298
p mux3_1x_8_0/mux3_dp_1x_5/a_33_7# result2 Vdd! 2 10 355 297
n mux3_1x_8_0/mux3_dp_1x_7/s0 mux3_1x_8_0/mux3_dp_1x_5/a_0_7# mux3_1x_8_0/mux3_dp_1x_5/a_7_7# 2 6 301 231
n adder_8_0/b_2_ mux3_1x_8_0/mux3_dp_1x_5/a_7_7# Gnd! 2 6 306 231
n adder_8_0/s_2_ Gnd! mux3_1x_8_0/mux3_dp_1x_5/a_20_7# 2 6 314 231
n mux3_1x_8_0/mux3_dp_1x_7/s0b mux3_1x_8_0/mux3_dp_1x_5/a_20_7# mux3_1x_8_0/mux3_dp_1x_5/a_0_7# 2 6 319 231
n mux3_1x_8_0/mux3_dp_1x_7/s1b mux3_1x_8_0/mux3_dp_1x_5/a_0_7# mux3_1x_8_0/mux3_dp_1x_5/a_33_7# 2 6 327 231
n mux3_1x_8_0/mux3_dp_1x_7/s1 mux3_1x_8_0/mux3_dp_1x_5/a_33_7# mux3_1x_8_0/mux3_dp_1x_5/a_41_7# 2 6 335 231
n less mux3_1x_8_0/mux3_dp_1x_5/a_41_7# Gnd! 2 6 340 231
n mux3_1x_8_0/mux3_dp_1x_5/a_33_7# Gnd! result2 2 7 358 236
p mux3_1x_8_0/mux3_dp_1x_7/s0 mux3_1x_8_0/mux3_dp_1x_4/a_0_74# mux3_1x_8_0/mux3_dp_1x_4/a_7_74# 2 9 301 408
p adder_8_0/s_3_ mux3_1x_8_0/mux3_dp_1x_4/a_7_74# Vdd! 2 9 306 408
p adder_8_0/b_3_ Vdd! mux3_1x_8_0/mux3_dp_1x_4/a_20_74# 2 9 314 408
p mux3_1x_8_0/mux3_dp_1x_7/s0b mux3_1x_8_0/mux3_dp_1x_4/a_20_74# mux3_1x_8_0/mux3_dp_1x_4/a_0_74# 2 9 319 408
p mux3_1x_8_0/mux3_dp_1x_7/s1 mux3_1x_8_0/mux3_dp_1x_4/a_0_74# mux3_1x_8_0/mux3_dp_1x_4/a_33_7# 2 9 327 408
p mux3_1x_8_0/mux3_dp_1x_7/s1b mux3_1x_8_0/mux3_dp_1x_4/a_33_7# mux3_1x_8_0/mux3_dp_1x_4/a_41_74# 2 9 335 408
p less mux3_1x_8_0/mux3_dp_1x_4/a_41_74# Vdd! 2 9 340 408
p mux3_1x_8_0/mux3_dp_1x_4/a_33_7# result3 Vdd! 2 10 355 407
n mux3_1x_8_0/mux3_dp_1x_7/s0 mux3_1x_8_0/mux3_dp_1x_4/a_0_7# mux3_1x_8_0/mux3_dp_1x_4/a_7_7# 2 6 301 341
n adder_8_0/b_3_ mux3_1x_8_0/mux3_dp_1x_4/a_7_7# Gnd! 2 6 306 341
n adder_8_0/s_3_ Gnd! mux3_1x_8_0/mux3_dp_1x_4/a_20_7# 2 6 314 341
n mux3_1x_8_0/mux3_dp_1x_7/s0b mux3_1x_8_0/mux3_dp_1x_4/a_20_7# mux3_1x_8_0/mux3_dp_1x_4/a_0_7# 2 6 319 341
n mux3_1x_8_0/mux3_dp_1x_7/s1b mux3_1x_8_0/mux3_dp_1x_4/a_0_7# mux3_1x_8_0/mux3_dp_1x_4/a_33_7# 2 6 327 341
n mux3_1x_8_0/mux3_dp_1x_7/s1 mux3_1x_8_0/mux3_dp_1x_4/a_33_7# mux3_1x_8_0/mux3_dp_1x_4/a_41_7# 2 6 335 341
n less mux3_1x_8_0/mux3_dp_1x_4/a_41_7# Gnd! 2 6 340 341
n mux3_1x_8_0/mux3_dp_1x_4/a_33_7# Gnd! result3 2 7 358 346
p mux3_1x_8_0/mux3_dp_1x_7/s0 mux3_1x_8_0/mux3_dp_1x_3/a_0_74# mux3_1x_8_0/mux3_dp_1x_3/a_7_74# 2 9 301 518
p adder_8_0/s_4_ mux3_1x_8_0/mux3_dp_1x_3/a_7_74# Vdd! 2 9 306 518
p adder_8_0/b_4_ Vdd! mux3_1x_8_0/mux3_dp_1x_3/a_20_74# 2 9 314 518
p mux3_1x_8_0/mux3_dp_1x_7/s0b mux3_1x_8_0/mux3_dp_1x_3/a_20_74# mux3_1x_8_0/mux3_dp_1x_3/a_0_74# 2 9 319 518
p mux3_1x_8_0/mux3_dp_1x_7/s1 mux3_1x_8_0/mux3_dp_1x_3/a_0_74# mux3_1x_8_0/mux3_dp_1x_3/a_33_7# 2 9 327 518
p mux3_1x_8_0/mux3_dp_1x_7/s1b mux3_1x_8_0/mux3_dp_1x_3/a_33_7# mux3_1x_8_0/mux3_dp_1x_3/a_41_74# 2 9 335 518
p less mux3_1x_8_0/mux3_dp_1x_3/a_41_74# Vdd! 2 9 340 518
p mux3_1x_8_0/mux3_dp_1x_3/a_33_7# result4 Vdd! 2 10 355 517
n mux3_1x_8_0/mux3_dp_1x_7/s0 mux3_1x_8_0/mux3_dp_1x_3/a_0_7# mux3_1x_8_0/mux3_dp_1x_3/a_7_7# 2 6 301 451
n adder_8_0/b_4_ mux3_1x_8_0/mux3_dp_1x_3/a_7_7# Gnd! 2 6 306 451
n adder_8_0/s_4_ Gnd! mux3_1x_8_0/mux3_dp_1x_3/a_20_7# 2 6 314 451
n mux3_1x_8_0/mux3_dp_1x_7/s0b mux3_1x_8_0/mux3_dp_1x_3/a_20_7# mux3_1x_8_0/mux3_dp_1x_3/a_0_7# 2 6 319 451
n mux3_1x_8_0/mux3_dp_1x_7/s1b mux3_1x_8_0/mux3_dp_1x_3/a_0_7# mux3_1x_8_0/mux3_dp_1x_3/a_33_7# 2 6 327 451
n mux3_1x_8_0/mux3_dp_1x_7/s1 mux3_1x_8_0/mux3_dp_1x_3/a_33_7# mux3_1x_8_0/mux3_dp_1x_3/a_41_7# 2 6 335 451
n less mux3_1x_8_0/mux3_dp_1x_3/a_41_7# Gnd! 2 6 340 451
n mux3_1x_8_0/mux3_dp_1x_3/a_33_7# Gnd! result4 2 7 358 456
p mux3_1x_8_0/mux3_dp_1x_7/s0 mux3_1x_8_0/mux3_dp_1x_2/a_0_74# mux3_1x_8_0/mux3_dp_1x_2/a_7_74# 2 9 301 628
p adder_8_0/s_5_ mux3_1x_8_0/mux3_dp_1x_2/a_7_74# Vdd! 2 9 306 628
p adder_8_0/b_5_ Vdd! mux3_1x_8_0/mux3_dp_1x_2/a_20_74# 2 9 314 628
p mux3_1x_8_0/mux3_dp_1x_7/s0b mux3_1x_8_0/mux3_dp_1x_2/a_20_74# mux3_1x_8_0/mux3_dp_1x_2/a_0_74# 2 9 319 628
p mux3_1x_8_0/mux3_dp_1x_7/s1 mux3_1x_8_0/mux3_dp_1x_2/a_0_74# mux3_1x_8_0/mux3_dp_1x_2/a_33_7# 2 9 327 628
p mux3_1x_8_0/mux3_dp_1x_7/s1b mux3_1x_8_0/mux3_dp_1x_2/a_33_7# mux3_1x_8_0/mux3_dp_1x_2/a_41_74# 2 9 335 628
p less mux3_1x_8_0/mux3_dp_1x_2/a_41_74# Vdd! 2 9 340 628
p mux3_1x_8_0/mux3_dp_1x_2/a_33_7# result5 Vdd! 2 10 355 627
n mux3_1x_8_0/mux3_dp_1x_7/s0 mux3_1x_8_0/mux3_dp_1x_2/a_0_7# mux3_1x_8_0/mux3_dp_1x_2/a_7_7# 2 6 301 561
n adder_8_0/b_5_ mux3_1x_8_0/mux3_dp_1x_2/a_7_7# Gnd! 2 6 306 561
n adder_8_0/s_5_ Gnd! mux3_1x_8_0/mux3_dp_1x_2/a_20_7# 2 6 314 561
n mux3_1x_8_0/mux3_dp_1x_7/s0b mux3_1x_8_0/mux3_dp_1x_2/a_20_7# mux3_1x_8_0/mux3_dp_1x_2/a_0_7# 2 6 319 561
n mux3_1x_8_0/mux3_dp_1x_7/s1b mux3_1x_8_0/mux3_dp_1x_2/a_0_7# mux3_1x_8_0/mux3_dp_1x_2/a_33_7# 2 6 327 561
n mux3_1x_8_0/mux3_dp_1x_7/s1 mux3_1x_8_0/mux3_dp_1x_2/a_33_7# mux3_1x_8_0/mux3_dp_1x_2/a_41_7# 2 6 335 561
n less mux3_1x_8_0/mux3_dp_1x_2/a_41_7# Gnd! 2 6 340 561
n mux3_1x_8_0/mux3_dp_1x_2/a_33_7# Gnd! result5 2 7 358 566
p mux3_1x_8_0/mux3_dp_1x_7/s0 mux3_1x_8_0/mux3_dp_1x_1/a_0_74# mux3_1x_8_0/mux3_dp_1x_1/a_7_74# 2 9 301 738
p adder_8_0/s_6_ mux3_1x_8_0/mux3_dp_1x_1/a_7_74# Vdd! 2 9 306 738
p adder_8_0/b_6_ Vdd! mux3_1x_8_0/mux3_dp_1x_1/a_20_74# 2 9 314 738
p mux3_1x_8_0/mux3_dp_1x_7/s0b mux3_1x_8_0/mux3_dp_1x_1/a_20_74# mux3_1x_8_0/mux3_dp_1x_1/a_0_74# 2 9 319 738
p mux3_1x_8_0/mux3_dp_1x_7/s1 mux3_1x_8_0/mux3_dp_1x_1/a_0_74# mux3_1x_8_0/mux3_dp_1x_1/a_33_7# 2 9 327 738
p mux3_1x_8_0/mux3_dp_1x_7/s1b mux3_1x_8_0/mux3_dp_1x_1/a_33_7# mux3_1x_8_0/mux3_dp_1x_1/a_41_74# 2 9 335 738
p less mux3_1x_8_0/mux3_dp_1x_1/a_41_74# Vdd! 2 9 340 738
p mux3_1x_8_0/mux3_dp_1x_1/a_33_7# result6 Vdd! 2 10 355 737
n mux3_1x_8_0/mux3_dp_1x_7/s0 mux3_1x_8_0/mux3_dp_1x_1/a_0_7# mux3_1x_8_0/mux3_dp_1x_1/a_7_7# 2 6 301 671
n adder_8_0/b_6_ mux3_1x_8_0/mux3_dp_1x_1/a_7_7# Gnd! 2 6 306 671
n adder_8_0/s_6_ Gnd! mux3_1x_8_0/mux3_dp_1x_1/a_20_7# 2 6 314 671
n mux3_1x_8_0/mux3_dp_1x_7/s0b mux3_1x_8_0/mux3_dp_1x_1/a_20_7# mux3_1x_8_0/mux3_dp_1x_1/a_0_7# 2 6 319 671
n mux3_1x_8_0/mux3_dp_1x_7/s1b mux3_1x_8_0/mux3_dp_1x_1/a_0_7# mux3_1x_8_0/mux3_dp_1x_1/a_33_7# 2 6 327 671
n mux3_1x_8_0/mux3_dp_1x_7/s1 mux3_1x_8_0/mux3_dp_1x_1/a_33_7# mux3_1x_8_0/mux3_dp_1x_1/a_41_7# 2 6 335 671
n less mux3_1x_8_0/mux3_dp_1x_1/a_41_7# Gnd! 2 6 340 671
n mux3_1x_8_0/mux3_dp_1x_1/a_33_7# Gnd! result6 2 7 358 676
p mux3_1x_8_0/mux3_dp_1x_7/s0 mux3_1x_8_0/mux3_dp_1x_0/a_0_74# mux3_1x_8_0/mux3_dp_1x_0/a_7_74# 2 9 301 848
p adder_8_0/s_7_ mux3_1x_8_0/mux3_dp_1x_0/a_7_74# Vdd! 2 9 306 848
p adder_8_0/b_7_ Vdd! mux3_1x_8_0/mux3_dp_1x_0/a_20_74# 2 9 314 848
p mux3_1x_8_0/mux3_dp_1x_7/s0b mux3_1x_8_0/mux3_dp_1x_0/a_20_74# mux3_1x_8_0/mux3_dp_1x_0/a_0_74# 2 9 319 848
p mux3_1x_8_0/mux3_dp_1x_7/s1 mux3_1x_8_0/mux3_dp_1x_0/a_0_74# mux3_1x_8_0/mux3_dp_1x_0/a_33_7# 2 9 327 848
p mux3_1x_8_0/mux3_dp_1x_7/s1b mux3_1x_8_0/mux3_dp_1x_0/a_33_7# mux3_1x_8_0/mux3_dp_1x_0/a_41_74# 2 9 335 848
p less mux3_1x_8_0/mux3_dp_1x_0/a_41_74# Vdd! 2 9 340 848
p mux3_1x_8_0/mux3_dp_1x_0/a_33_7# result7 Vdd! 2 10 355 847
n mux3_1x_8_0/mux3_dp_1x_7/s0 mux3_1x_8_0/mux3_dp_1x_0/a_0_7# mux3_1x_8_0/mux3_dp_1x_0/a_7_7# 2 6 301 781
n adder_8_0/b_7_ mux3_1x_8_0/mux3_dp_1x_0/a_7_7# Gnd! 2 6 306 781
n adder_8_0/s_7_ Gnd! mux3_1x_8_0/mux3_dp_1x_0/a_20_7# 2 6 314 781
n mux3_1x_8_0/mux3_dp_1x_7/s0b mux3_1x_8_0/mux3_dp_1x_0/a_20_7# mux3_1x_8_0/mux3_dp_1x_0/a_0_7# 2 6 319 781
n mux3_1x_8_0/mux3_dp_1x_7/s1b mux3_1x_8_0/mux3_dp_1x_0/a_0_7# mux3_1x_8_0/mux3_dp_1x_0/a_33_7# 2 6 327 781
n mux3_1x_8_0/mux3_dp_1x_7/s1 mux3_1x_8_0/mux3_dp_1x_0/a_33_7# mux3_1x_8_0/mux3_dp_1x_0/a_41_7# 2 6 335 781
n less mux3_1x_8_0/mux3_dp_1x_0/a_41_7# Gnd! 2 6 340 781
n mux3_1x_8_0/mux3_dp_1x_0/a_33_7# Gnd! result7 2 7 358 786
p op1 Vdd! mux3_1x_8_0/mux3_dp_1x_7/s1b 2 37 333 930
p mux3_1x_8_0/mux3_dp_1x_7/s1b Vdd! mux3_1x_8_0/mux3_dp_1x_7/s1 2 37 349 930
n op1 Gnd! mux3_1x_8_0/mux3_dp_1x_7/s1b 2 27 333 891
n mux3_1x_8_0/mux3_dp_1x_7/s1b Gnd! mux3_1x_8_0/mux3_dp_1x_7/s1 2 27 349 891
p op0 Vdd! mux3_1x_8_0/mux3_dp_1x_7/s0b 2 37 301 930
p mux3_1x_8_0/mux3_dp_1x_7/s0b Vdd! mux3_1x_8_0/mux3_dp_1x_7/s0 2 37 317 930
n op0 Gnd! mux3_1x_8_0/mux3_dp_1x_7/s0b 2 27 301 891
n mux3_1x_8_0/mux3_dp_1x_7/s0b Gnd! mux3_1x_8_0/mux3_dp_1x_7/s0 2 27 317 891
p a0 adder_8_0/fulladder_7/a_n2_65# Vdd! 2 16 173 69
p muxy7 Vdd! adder_8_0/fulladder_7/a_n2_65# 2 16 181 69
p op2 adder_8_0/fulladder_7/a_n2_65# adder_8_0/fulladder_7/a_21_7# 2 16 189 69
p muxy7 adder_8_0/fulladder_7/a_21_7# adder_8_0/fulladder_7/a_29_65# 2 16 197 69
p a0 adder_8_0/fulladder_7/a_29_65# Vdd! 2 16 205 69
p a0 Vdd! adder_8_0/fulladder_7/a_45_65# 2 16 213 69
p muxy7 adder_8_0/fulladder_7/a_45_65# Vdd! 2 16 221 69
p op2 Vdd! adder_8_0/fulladder_7/a_45_65# 2 16 229 69
p adder_8_0/fulladder_7/a_21_7# adder_8_0/fulladder_7/a_45_65# adder_8_0/fulladder_7/a_69_7# 2 16 237 69
p op2 adder_8_0/fulladder_7/a_69_7# adder_8_0/fulladder_7/a_77_65# 2 16 245 69
p muxy7 adder_8_0/fulladder_7/a_77_65# adder_8_0/fulladder_7/a_85_65# 2 16 253 69
p a0 adder_8_0/fulladder_7/a_85_65# Vdd! 2 16 261 69
p adder_8_0/fulladder_7/a_69_7# Vdd! adder_8_0/s_0_ 2 16 269 69
p adder_8_0/fulladder_7/a_21_7# Vdd! adder_8_0/c_1_ 2 16 285 69
n a0 adder_8_0/fulladder_7/a_n2_7# Gnd! 2 8 173 11
n muxy7 Gnd! adder_8_0/fulladder_7/a_n2_7# 2 8 181 11
n op2 adder_8_0/fulladder_7/a_n2_7# adder_8_0/fulladder_7/a_21_7# 2 8 189 11
n muxy7 adder_8_0/fulladder_7/a_21_7# adder_8_0/fulladder_7/a_29_7# 2 8 197 11
n a0 adder_8_0/fulladder_7/a_29_7# Gnd! 2 8 205 11
n a0 Gnd! adder_8_0/fulladder_7/a_45_7# 2 8 213 11
n muxy7 adder_8_0/fulladder_7/a_45_7# Gnd! 2 8 221 11
n op2 Gnd! adder_8_0/fulladder_7/a_45_7# 2 8 229 11
n adder_8_0/fulladder_7/a_21_7# adder_8_0/fulladder_7/a_45_7# adder_8_0/fulladder_7/a_69_7# 2 8 237 11
n op2 adder_8_0/fulladder_7/a_69_7# adder_8_0/fulladder_7/a_77_7# 2 8 245 11
n muxy7 adder_8_0/fulladder_7/a_77_7# adder_8_0/fulladder_7/a_85_7# 2 8 253 11
n a0 adder_8_0/fulladder_7/a_85_7# Gnd! 2 8 261 11
n adder_8_0/fulladder_7/a_69_7# Gnd! adder_8_0/s_0_ 2 8 269 11
n adder_8_0/fulladder_7/a_21_7# Gnd! adder_8_0/c_1_ 2 8 285 11
p a1 adder_8_0/fulladder_6/a_n2_65# Vdd! 2 16 173 179
p adder_8_0/b_1_ Vdd! adder_8_0/fulladder_6/a_n2_65# 2 16 181 179
p adder_8_0/c_1_ adder_8_0/fulladder_6/a_n2_65# adder_8_0/fulladder_6/a_21_7# 2 16 189 179
p adder_8_0/b_1_ adder_8_0/fulladder_6/a_21_7# adder_8_0/fulladder_6/a_29_65# 2 16 197 179
p a1 adder_8_0/fulladder_6/a_29_65# Vdd! 2 16 205 179
p a1 Vdd! adder_8_0/fulladder_6/a_45_65# 2 16 213 179
p adder_8_0/b_1_ adder_8_0/fulladder_6/a_45_65# Vdd! 2 16 221 179
p adder_8_0/c_1_ Vdd! adder_8_0/fulladder_6/a_45_65# 2 16 229 179
p adder_8_0/fulladder_6/a_21_7# adder_8_0/fulladder_6/a_45_65# adder_8_0/fulladder_6/a_69_7# 2 16 237 179
p adder_8_0/c_1_ adder_8_0/fulladder_6/a_69_7# adder_8_0/fulladder_6/a_77_65# 2 16 245 179
p adder_8_0/b_1_ adder_8_0/fulladder_6/a_77_65# adder_8_0/fulladder_6/a_85_65# 2 16 253 179
p a1 adder_8_0/fulladder_6/a_85_65# Vdd! 2 16 261 179
p adder_8_0/fulladder_6/a_69_7# Vdd! adder_8_0/s_1_ 2 16 269 179
p adder_8_0/fulladder_6/a_21_7# Vdd! adder_8_0/c_2_ 2 16 285 179
n a1 adder_8_0/fulladder_6/a_n2_7# Gnd! 2 8 173 121
n adder_8_0/b_1_ Gnd! adder_8_0/fulladder_6/a_n2_7# 2 8 181 121
n adder_8_0/c_1_ adder_8_0/fulladder_6/a_n2_7# adder_8_0/fulladder_6/a_21_7# 2 8 189 121
n adder_8_0/b_1_ adder_8_0/fulladder_6/a_21_7# adder_8_0/fulladder_6/a_29_7# 2 8 197 121
n a1 adder_8_0/fulladder_6/a_29_7# Gnd! 2 8 205 121
n a1 Gnd! adder_8_0/fulladder_6/a_45_7# 2 8 213 121
n adder_8_0/b_1_ adder_8_0/fulladder_6/a_45_7# Gnd! 2 8 221 121
n adder_8_0/c_1_ Gnd! adder_8_0/fulladder_6/a_45_7# 2 8 229 121
n adder_8_0/fulladder_6/a_21_7# adder_8_0/fulladder_6/a_45_7# adder_8_0/fulladder_6/a_69_7# 2 8 237 121
n adder_8_0/c_1_ adder_8_0/fulladder_6/a_69_7# adder_8_0/fulladder_6/a_77_7# 2 8 245 121
n adder_8_0/b_1_ adder_8_0/fulladder_6/a_77_7# adder_8_0/fulladder_6/a_85_7# 2 8 253 121
n a1 adder_8_0/fulladder_6/a_85_7# Gnd! 2 8 261 121
n adder_8_0/fulladder_6/a_69_7# Gnd! adder_8_0/s_1_ 2 8 269 121
n adder_8_0/fulladder_6/a_21_7# Gnd! adder_8_0/c_2_ 2 8 285 121
p a2 adder_8_0/fulladder_5/a_n2_65# Vdd! 2 16 173 289
p adder_8_0/b_2_ Vdd! adder_8_0/fulladder_5/a_n2_65# 2 16 181 289
p adder_8_0/c_2_ adder_8_0/fulladder_5/a_n2_65# adder_8_0/fulladder_5/a_21_7# 2 16 189 289
p adder_8_0/b_2_ adder_8_0/fulladder_5/a_21_7# adder_8_0/fulladder_5/a_29_65# 2 16 197 289
p a2 adder_8_0/fulladder_5/a_29_65# Vdd! 2 16 205 289
p a2 Vdd! adder_8_0/fulladder_5/a_45_65# 2 16 213 289
p adder_8_0/b_2_ adder_8_0/fulladder_5/a_45_65# Vdd! 2 16 221 289
p adder_8_0/c_2_ Vdd! adder_8_0/fulladder_5/a_45_65# 2 16 229 289
p adder_8_0/fulladder_5/a_21_7# adder_8_0/fulladder_5/a_45_65# adder_8_0/fulladder_5/a_69_7# 2 16 237 289
p adder_8_0/c_2_ adder_8_0/fulladder_5/a_69_7# adder_8_0/fulladder_5/a_77_65# 2 16 245 289
p adder_8_0/b_2_ adder_8_0/fulladder_5/a_77_65# adder_8_0/fulladder_5/a_85_65# 2 16 253 289
p a2 adder_8_0/fulladder_5/a_85_65# Vdd! 2 16 261 289
p adder_8_0/fulladder_5/a_69_7# Vdd! adder_8_0/s_2_ 2 16 269 289
p adder_8_0/fulladder_5/a_21_7# Vdd! adder_8_0/c_3_ 2 16 285 289
n a2 adder_8_0/fulladder_5/a_n2_7# Gnd! 2 8 173 231
n adder_8_0/b_2_ Gnd! adder_8_0/fulladder_5/a_n2_7# 2 8 181 231
n adder_8_0/c_2_ adder_8_0/fulladder_5/a_n2_7# adder_8_0/fulladder_5/a_21_7# 2 8 189 231
n adder_8_0/b_2_ adder_8_0/fulladder_5/a_21_7# adder_8_0/fulladder_5/a_29_7# 2 8 197 231
n a2 adder_8_0/fulladder_5/a_29_7# Gnd! 2 8 205 231
n a2 Gnd! adder_8_0/fulladder_5/a_45_7# 2 8 213 231
n adder_8_0/b_2_ adder_8_0/fulladder_5/a_45_7# Gnd! 2 8 221 231
n adder_8_0/c_2_ Gnd! adder_8_0/fulladder_5/a_45_7# 2 8 229 231
n adder_8_0/fulladder_5/a_21_7# adder_8_0/fulladder_5/a_45_7# adder_8_0/fulladder_5/a_69_7# 2 8 237 231
n adder_8_0/c_2_ adder_8_0/fulladder_5/a_69_7# adder_8_0/fulladder_5/a_77_7# 2 8 245 231
n adder_8_0/b_2_ adder_8_0/fulladder_5/a_77_7# adder_8_0/fulladder_5/a_85_7# 2 8 253 231
n a2 adder_8_0/fulladder_5/a_85_7# Gnd! 2 8 261 231
n adder_8_0/fulladder_5/a_69_7# Gnd! adder_8_0/s_2_ 2 8 269 231
n adder_8_0/fulladder_5/a_21_7# Gnd! adder_8_0/c_3_ 2 8 285 231
p a3 adder_8_0/fulladder_4/a_n2_65# Vdd! 2 16 173 399
p adder_8_0/b_3_ Vdd! adder_8_0/fulladder_4/a_n2_65# 2 16 181 399
p adder_8_0/c_3_ adder_8_0/fulladder_4/a_n2_65# adder_8_0/fulladder_4/a_21_7# 2 16 189 399
p adder_8_0/b_3_ adder_8_0/fulladder_4/a_21_7# adder_8_0/fulladder_4/a_29_65# 2 16 197 399
p a3 adder_8_0/fulladder_4/a_29_65# Vdd! 2 16 205 399
p a3 Vdd! adder_8_0/fulladder_4/a_45_65# 2 16 213 399
p adder_8_0/b_3_ adder_8_0/fulladder_4/a_45_65# Vdd! 2 16 221 399
p adder_8_0/c_3_ Vdd! adder_8_0/fulladder_4/a_45_65# 2 16 229 399
p adder_8_0/fulladder_4/a_21_7# adder_8_0/fulladder_4/a_45_65# adder_8_0/fulladder_4/a_69_7# 2 16 237 399
p adder_8_0/c_3_ adder_8_0/fulladder_4/a_69_7# adder_8_0/fulladder_4/a_77_65# 2 16 245 399
p adder_8_0/b_3_ adder_8_0/fulladder_4/a_77_65# adder_8_0/fulladder_4/a_85_65# 2 16 253 399
p a3 adder_8_0/fulladder_4/a_85_65# Vdd! 2 16 261 399
p adder_8_0/fulladder_4/a_69_7# Vdd! adder_8_0/s_3_ 2 16 269 399
p adder_8_0/fulladder_4/a_21_7# Vdd! adder_8_0/c_4_ 2 16 285 399
n a3 adder_8_0/fulladder_4/a_n2_7# Gnd! 2 8 173 341
n adder_8_0/b_3_ Gnd! adder_8_0/fulladder_4/a_n2_7# 2 8 181 341
n adder_8_0/c_3_ adder_8_0/fulladder_4/a_n2_7# adder_8_0/fulladder_4/a_21_7# 2 8 189 341
n adder_8_0/b_3_ adder_8_0/fulladder_4/a_21_7# adder_8_0/fulladder_4/a_29_7# 2 8 197 341
n a3 adder_8_0/fulladder_4/a_29_7# Gnd! 2 8 205 341
n a3 Gnd! adder_8_0/fulladder_4/a_45_7# 2 8 213 341
n adder_8_0/b_3_ adder_8_0/fulladder_4/a_45_7# Gnd! 2 8 221 341
n adder_8_0/c_3_ Gnd! adder_8_0/fulladder_4/a_45_7# 2 8 229 341
n adder_8_0/fulladder_4/a_21_7# adder_8_0/fulladder_4/a_45_7# adder_8_0/fulladder_4/a_69_7# 2 8 237 341
n adder_8_0/c_3_ adder_8_0/fulladder_4/a_69_7# adder_8_0/fulladder_4/a_77_7# 2 8 245 341
n adder_8_0/b_3_ adder_8_0/fulladder_4/a_77_7# adder_8_0/fulladder_4/a_85_7# 2 8 253 341
n a3 adder_8_0/fulladder_4/a_85_7# Gnd! 2 8 261 341
n adder_8_0/fulladder_4/a_69_7# Gnd! adder_8_0/s_3_ 2 8 269 341
n adder_8_0/fulladder_4/a_21_7# Gnd! adder_8_0/c_4_ 2 8 285 341
p a4 adder_8_0/fulladder_3/a_n2_65# Vdd! 2 16 173 509
p adder_8_0/b_4_ Vdd! adder_8_0/fulladder_3/a_n2_65# 2 16 181 509
p adder_8_0/c_4_ adder_8_0/fulladder_3/a_n2_65# adder_8_0/fulladder_3/a_21_7# 2 16 189 509
p adder_8_0/b_4_ adder_8_0/fulladder_3/a_21_7# adder_8_0/fulladder_3/a_29_65# 2 16 197 509
p a4 adder_8_0/fulladder_3/a_29_65# Vdd! 2 16 205 509
p a4 Vdd! adder_8_0/fulladder_3/a_45_65# 2 16 213 509
p adder_8_0/b_4_ adder_8_0/fulladder_3/a_45_65# Vdd! 2 16 221 509
p adder_8_0/c_4_ Vdd! adder_8_0/fulladder_3/a_45_65# 2 16 229 509
p adder_8_0/fulladder_3/a_21_7# adder_8_0/fulladder_3/a_45_65# adder_8_0/fulladder_3/a_69_7# 2 16 237 509
p adder_8_0/c_4_ adder_8_0/fulladder_3/a_69_7# adder_8_0/fulladder_3/a_77_65# 2 16 245 509
p adder_8_0/b_4_ adder_8_0/fulladder_3/a_77_65# adder_8_0/fulladder_3/a_85_65# 2 16 253 509
p a4 adder_8_0/fulladder_3/a_85_65# Vdd! 2 16 261 509
p adder_8_0/fulladder_3/a_69_7# Vdd! adder_8_0/s_4_ 2 16 269 509
p adder_8_0/fulladder_3/a_21_7# Vdd! adder_8_0/c_5_ 2 16 285 509
n a4 adder_8_0/fulladder_3/a_n2_7# Gnd! 2 8 173 451
n adder_8_0/b_4_ Gnd! adder_8_0/fulladder_3/a_n2_7# 2 8 181 451
n adder_8_0/c_4_ adder_8_0/fulladder_3/a_n2_7# adder_8_0/fulladder_3/a_21_7# 2 8 189 451
n adder_8_0/b_4_ adder_8_0/fulladder_3/a_21_7# adder_8_0/fulladder_3/a_29_7# 2 8 197 451
n a4 adder_8_0/fulladder_3/a_29_7# Gnd! 2 8 205 451
n a4 Gnd! adder_8_0/fulladder_3/a_45_7# 2 8 213 451
n adder_8_0/b_4_ adder_8_0/fulladder_3/a_45_7# Gnd! 2 8 221 451
n adder_8_0/c_4_ Gnd! adder_8_0/fulladder_3/a_45_7# 2 8 229 451
n adder_8_0/fulladder_3/a_21_7# adder_8_0/fulladder_3/a_45_7# adder_8_0/fulladder_3/a_69_7# 2 8 237 451
n adder_8_0/c_4_ adder_8_0/fulladder_3/a_69_7# adder_8_0/fulladder_3/a_77_7# 2 8 245 451
n adder_8_0/b_4_ adder_8_0/fulladder_3/a_77_7# adder_8_0/fulladder_3/a_85_7# 2 8 253 451
n a4 adder_8_0/fulladder_3/a_85_7# Gnd! 2 8 261 451
n adder_8_0/fulladder_3/a_69_7# Gnd! adder_8_0/s_4_ 2 8 269 451
n adder_8_0/fulladder_3/a_21_7# Gnd! adder_8_0/c_5_ 2 8 285 451
p a5 adder_8_0/fulladder_2/a_n2_65# Vdd! 2 16 173 619
p adder_8_0/b_5_ Vdd! adder_8_0/fulladder_2/a_n2_65# 2 16 181 619
p adder_8_0/c_5_ adder_8_0/fulladder_2/a_n2_65# adder_8_0/fulladder_2/a_21_7# 2 16 189 619
p adder_8_0/b_5_ adder_8_0/fulladder_2/a_21_7# adder_8_0/fulladder_2/a_29_65# 2 16 197 619
p a5 adder_8_0/fulladder_2/a_29_65# Vdd! 2 16 205 619
p a5 Vdd! adder_8_0/fulladder_2/a_45_65# 2 16 213 619
p adder_8_0/b_5_ adder_8_0/fulladder_2/a_45_65# Vdd! 2 16 221 619
p adder_8_0/c_5_ Vdd! adder_8_0/fulladder_2/a_45_65# 2 16 229 619
p adder_8_0/fulladder_2/a_21_7# adder_8_0/fulladder_2/a_45_65# adder_8_0/fulladder_2/a_69_7# 2 16 237 619
p adder_8_0/c_5_ adder_8_0/fulladder_2/a_69_7# adder_8_0/fulladder_2/a_77_65# 2 16 245 619
p adder_8_0/b_5_ adder_8_0/fulladder_2/a_77_65# adder_8_0/fulladder_2/a_85_65# 2 16 253 619
p a5 adder_8_0/fulladder_2/a_85_65# Vdd! 2 16 261 619
p adder_8_0/fulladder_2/a_69_7# Vdd! adder_8_0/s_5_ 2 16 269 619
p adder_8_0/fulladder_2/a_21_7# Vdd! adder_8_0/c_6_ 2 16 285 619
n a5 adder_8_0/fulladder_2/a_n2_7# Gnd! 2 8 173 561
n adder_8_0/b_5_ Gnd! adder_8_0/fulladder_2/a_n2_7# 2 8 181 561
n adder_8_0/c_5_ adder_8_0/fulladder_2/a_n2_7# adder_8_0/fulladder_2/a_21_7# 2 8 189 561
n adder_8_0/b_5_ adder_8_0/fulladder_2/a_21_7# adder_8_0/fulladder_2/a_29_7# 2 8 197 561
n a5 adder_8_0/fulladder_2/a_29_7# Gnd! 2 8 205 561
n a5 Gnd! adder_8_0/fulladder_2/a_45_7# 2 8 213 561
n adder_8_0/b_5_ adder_8_0/fulladder_2/a_45_7# Gnd! 2 8 221 561
n adder_8_0/c_5_ Gnd! adder_8_0/fulladder_2/a_45_7# 2 8 229 561
n adder_8_0/fulladder_2/a_21_7# adder_8_0/fulladder_2/a_45_7# adder_8_0/fulladder_2/a_69_7# 2 8 237 561
n adder_8_0/c_5_ adder_8_0/fulladder_2/a_69_7# adder_8_0/fulladder_2/a_77_7# 2 8 245 561
n adder_8_0/b_5_ adder_8_0/fulladder_2/a_77_7# adder_8_0/fulladder_2/a_85_7# 2 8 253 561
n a5 adder_8_0/fulladder_2/a_85_7# Gnd! 2 8 261 561
n adder_8_0/fulladder_2/a_69_7# Gnd! adder_8_0/s_5_ 2 8 269 561
n adder_8_0/fulladder_2/a_21_7# Gnd! adder_8_0/c_6_ 2 8 285 561
p a6 adder_8_0/fulladder_1/a_n2_65# Vdd! 2 16 173 729
p adder_8_0/b_6_ Vdd! adder_8_0/fulladder_1/a_n2_65# 2 16 181 729
p adder_8_0/c_6_ adder_8_0/fulladder_1/a_n2_65# adder_8_0/fulladder_1/a_21_7# 2 16 189 729
p adder_8_0/b_6_ adder_8_0/fulladder_1/a_21_7# adder_8_0/fulladder_1/a_29_65# 2 16 197 729
p a6 adder_8_0/fulladder_1/a_29_65# Vdd! 2 16 205 729
p a6 Vdd! adder_8_0/fulladder_1/a_45_65# 2 16 213 729
p adder_8_0/b_6_ adder_8_0/fulladder_1/a_45_65# Vdd! 2 16 221 729
p adder_8_0/c_6_ Vdd! adder_8_0/fulladder_1/a_45_65# 2 16 229 729
p adder_8_0/fulladder_1/a_21_7# adder_8_0/fulladder_1/a_45_65# adder_8_0/fulladder_1/a_69_7# 2 16 237 729
p adder_8_0/c_6_ adder_8_0/fulladder_1/a_69_7# adder_8_0/fulladder_1/a_77_65# 2 16 245 729
p adder_8_0/b_6_ adder_8_0/fulladder_1/a_77_65# adder_8_0/fulladder_1/a_85_65# 2 16 253 729
p a6 adder_8_0/fulladder_1/a_85_65# Vdd! 2 16 261 729
p adder_8_0/fulladder_1/a_69_7# Vdd! adder_8_0/s_6_ 2 16 269 729
p adder_8_0/fulladder_1/a_21_7# Vdd! adder_8_0/c_7_ 2 16 285 729
n a6 adder_8_0/fulladder_1/a_n2_7# Gnd! 2 8 173 671
n adder_8_0/b_6_ Gnd! adder_8_0/fulladder_1/a_n2_7# 2 8 181 671
n adder_8_0/c_6_ adder_8_0/fulladder_1/a_n2_7# adder_8_0/fulladder_1/a_21_7# 2 8 189 671
n adder_8_0/b_6_ adder_8_0/fulladder_1/a_21_7# adder_8_0/fulladder_1/a_29_7# 2 8 197 671
n a6 adder_8_0/fulladder_1/a_29_7# Gnd! 2 8 205 671
n a6 Gnd! adder_8_0/fulladder_1/a_45_7# 2 8 213 671
n adder_8_0/b_6_ adder_8_0/fulladder_1/a_45_7# Gnd! 2 8 221 671
n adder_8_0/c_6_ Gnd! adder_8_0/fulladder_1/a_45_7# 2 8 229 671
n adder_8_0/fulladder_1/a_21_7# adder_8_0/fulladder_1/a_45_7# adder_8_0/fulladder_1/a_69_7# 2 8 237 671
n adder_8_0/c_6_ adder_8_0/fulladder_1/a_69_7# adder_8_0/fulladder_1/a_77_7# 2 8 245 671
n adder_8_0/b_6_ adder_8_0/fulladder_1/a_77_7# adder_8_0/fulladder_1/a_85_7# 2 8 253 671
n a6 adder_8_0/fulladder_1/a_85_7# Gnd! 2 8 261 671
n adder_8_0/fulladder_1/a_69_7# Gnd! adder_8_0/s_6_ 2 8 269 671
n adder_8_0/fulladder_1/a_21_7# Gnd! adder_8_0/c_7_ 2 8 285 671
p a7 adder_8_0/fulladder_0/a_n2_65# Vdd! 2 16 173 839
p adder_8_0/b_7_ Vdd! adder_8_0/fulladder_0/a_n2_65# 2 16 181 839
p adder_8_0/c_7_ adder_8_0/fulladder_0/a_n2_65# adder_8_0/fulladder_0/a_21_7# 2 16 189 839
p adder_8_0/b_7_ adder_8_0/fulladder_0/a_21_7# adder_8_0/fulladder_0/a_29_65# 2 16 197 839
p a7 adder_8_0/fulladder_0/a_29_65# Vdd! 2 16 205 839
p a7 Vdd! adder_8_0/fulladder_0/a_45_65# 2 16 213 839
p adder_8_0/b_7_ adder_8_0/fulladder_0/a_45_65# Vdd! 2 16 221 839
p adder_8_0/c_7_ Vdd! adder_8_0/fulladder_0/a_45_65# 2 16 229 839
p adder_8_0/fulladder_0/a_21_7# adder_8_0/fulladder_0/a_45_65# adder_8_0/fulladder_0/a_69_7# 2 16 237 839
p adder_8_0/c_7_ adder_8_0/fulladder_0/a_69_7# adder_8_0/fulladder_0/a_77_65# 2 16 245 839
p adder_8_0/b_7_ adder_8_0/fulladder_0/a_77_65# adder_8_0/fulladder_0/a_85_65# 2 16 253 839
p a7 adder_8_0/fulladder_0/a_85_65# Vdd! 2 16 261 839
p adder_8_0/fulladder_0/a_69_7# Vdd! adder_8_0/s_7_ 2 16 269 839
p adder_8_0/fulladder_0/a_21_7# Vdd! cout_adder_7 2 16 285 839
n a7 adder_8_0/fulladder_0/a_n2_7# Gnd! 2 8 173 781
n adder_8_0/b_7_ Gnd! adder_8_0/fulladder_0/a_n2_7# 2 8 181 781
n adder_8_0/c_7_ adder_8_0/fulladder_0/a_n2_7# adder_8_0/fulladder_0/a_21_7# 2 8 189 781
n adder_8_0/b_7_ adder_8_0/fulladder_0/a_21_7# adder_8_0/fulladder_0/a_29_7# 2 8 197 781
n a7 adder_8_0/fulladder_0/a_29_7# Gnd! 2 8 205 781
n a7 Gnd! adder_8_0/fulladder_0/a_45_7# 2 8 213 781
n adder_8_0/b_7_ adder_8_0/fulladder_0/a_45_7# Gnd! 2 8 221 781
n adder_8_0/c_7_ Gnd! adder_8_0/fulladder_0/a_45_7# 2 8 229 781
n adder_8_0/fulladder_0/a_21_7# adder_8_0/fulladder_0/a_45_7# adder_8_0/fulladder_0/a_69_7# 2 8 237 781
n adder_8_0/c_7_ adder_8_0/fulladder_0/a_69_7# adder_8_0/fulladder_0/a_77_7# 2 8 245 781
n adder_8_0/b_7_ adder_8_0/fulladder_0/a_77_7# adder_8_0/fulladder_0/a_85_7# 2 8 253 781
n a7 adder_8_0/fulladder_0/a_85_7# Gnd! 2 8 261 781
n adder_8_0/fulladder_0/a_69_7# Gnd! adder_8_0/s_7_ 2 8 269 781
n adder_8_0/fulladder_0/a_21_7# Gnd! cout_adder_7 2 8 285 781
p b0 mux4_8_10space_0/mux4_dp_1x_0[0]/a_6_74# mux4_8_10space_0/mux4_dp_1x_0[0]/a_13_74# 2 9 75 78
p op6 mux4_8_10space_0/mux4_dp_1x_0[0]/a_13_74# Vdd! 2 9 80 78
p op5 Vdd! mux4_8_10space_0/mux4_dp_1x_0[0]/a_26_74# 2 9 88 78
p inv_1x_8_1/inv_1x_7/y mux4_8_10space_0/mux4_dp_1x_0[0]/a_26_74# mux4_8_10space_0/mux4_dp_1x_0[0]/a_6_74# 2 9 93 78
p a0 mux4_8_10space_0/mux4_dp_1x_0[0]/a_6_74# mux4_8_10space_0/mux4_dp_1x_0[0]/a_39_7# 2 9 101 78
p inv_1x_8_0/inv_1x_7/y mux4_8_10space_0/mux4_dp_1x_0[0]/a_39_7# mux4_8_10space_0/mux4_dp_1x_0[0]/a_47_74# 2 9 109 78
p b0 mux4_8_10space_0/mux4_dp_1x_0[0]/a_47_74# mux4_8_10space_0/mux4_dp_1x_0[0]/a_55_74# 2 9 117 78
p op4 mux4_8_10space_0/mux4_dp_1x_0[0]/a_55_74# Vdd! 2 9 122 78
p op3 Vdd! mux4_8_10space_0/mux4_dp_1x_0[0]/a_68_74# 2 9 130 78
p inv_1x_8_1/inv_1x_7/y mux4_8_10space_0/mux4_dp_1x_0[0]/a_68_74# mux4_8_10space_0/mux4_dp_1x_0[0]/a_47_74# 2 9 135 78
p mux4_8_10space_0/mux4_dp_1x_0[0]/a_39_7# Vdd! muxy7 2 10 157 77
n inv_1x_8_1/inv_1x_7/y mux4_8_10space_0/mux4_dp_1x_0[0]/a_6_7# mux4_8_10space_0/mux4_dp_1x_0[0]/a_13_7# 2 6 75 11
n op6 mux4_8_10space_0/mux4_dp_1x_0[0]/a_13_7# Gnd! 2 6 80 11
n op5 Gnd! mux4_8_10space_0/mux4_dp_1x_0[0]/a_26_7# 2 6 88 11
n b0 mux4_8_10space_0/mux4_dp_1x_0[0]/a_26_7# mux4_8_10space_0/mux4_dp_1x_0[0]/a_6_7# 2 6 93 11
n inv_1x_8_0/inv_1x_7/y mux4_8_10space_0/mux4_dp_1x_0[0]/a_6_7# mux4_8_10space_0/mux4_dp_1x_0[0]/a_39_7# 2 6 101 11
n a0 mux4_8_10space_0/mux4_dp_1x_0[0]/a_39_7# mux4_8_10space_0/mux4_dp_1x_0[0]/a_47_7# 2 6 109 11
n inv_1x_8_1/inv_1x_7/y mux4_8_10space_0/mux4_dp_1x_0[0]/a_47_7# mux4_8_10space_0/mux4_dp_1x_0[0]/a_55_7# 2 6 117 11
n op4 mux4_8_10space_0/mux4_dp_1x_0[0]/a_55_7# Gnd! 2 6 122 11
n op3 Gnd! mux4_8_10space_0/mux4_dp_1x_0[0]/a_68_7# 2 6 130 11
n b0 mux4_8_10space_0/mux4_dp_1x_0[0]/a_68_7# mux4_8_10space_0/mux4_dp_1x_0[0]/a_47_7# 2 6 135 11
n mux4_8_10space_0/mux4_dp_1x_0[0]/a_39_7# Gnd! muxy7 2 7 157 11
p b1 mux4_8_10space_0/mux4_dp_1x_0[1]/a_6_74# mux4_8_10space_0/mux4_dp_1x_0[1]/a_13_74# 2 9 75 188
p op6 mux4_8_10space_0/mux4_dp_1x_0[1]/a_13_74# Vdd! 2 9 80 188
p op5 Vdd! mux4_8_10space_0/mux4_dp_1x_0[1]/a_26_74# 2 9 88 188
p inv_1x_8_1/inv_1x_6/y mux4_8_10space_0/mux4_dp_1x_0[1]/a_26_74# mux4_8_10space_0/mux4_dp_1x_0[1]/a_6_74# 2 9 93 188
p a1 mux4_8_10space_0/mux4_dp_1x_0[1]/a_6_74# mux4_8_10space_0/mux4_dp_1x_0[1]/a_39_7# 2 9 101 188
p inv_1x_8_0/inv_1x_6/y mux4_8_10space_0/mux4_dp_1x_0[1]/a_39_7# mux4_8_10space_0/mux4_dp_1x_0[1]/a_47_74# 2 9 109 188
p b1 mux4_8_10space_0/mux4_dp_1x_0[1]/a_47_74# mux4_8_10space_0/mux4_dp_1x_0[1]/a_55_74# 2 9 117 188
p op4 mux4_8_10space_0/mux4_dp_1x_0[1]/a_55_74# Vdd! 2 9 122 188
p op3 Vdd! mux4_8_10space_0/mux4_dp_1x_0[1]/a_68_74# 2 9 130 188
p inv_1x_8_1/inv_1x_6/y mux4_8_10space_0/mux4_dp_1x_0[1]/a_68_74# mux4_8_10space_0/mux4_dp_1x_0[1]/a_47_74# 2 9 135 188
p mux4_8_10space_0/mux4_dp_1x_0[1]/a_39_7# Vdd! adder_8_0/b_1_ 2 10 157 187
n inv_1x_8_1/inv_1x_6/y mux4_8_10space_0/mux4_dp_1x_0[1]/a_6_7# mux4_8_10space_0/mux4_dp_1x_0[1]/a_13_7# 2 6 75 121
n op6 mux4_8_10space_0/mux4_dp_1x_0[1]/a_13_7# Gnd! 2 6 80 121
n op5 Gnd! mux4_8_10space_0/mux4_dp_1x_0[1]/a_26_7# 2 6 88 121
n b1 mux4_8_10space_0/mux4_dp_1x_0[1]/a_26_7# mux4_8_10space_0/mux4_dp_1x_0[1]/a_6_7# 2 6 93 121
n inv_1x_8_0/inv_1x_6/y mux4_8_10space_0/mux4_dp_1x_0[1]/a_6_7# mux4_8_10space_0/mux4_dp_1x_0[1]/a_39_7# 2 6 101 121
n a1 mux4_8_10space_0/mux4_dp_1x_0[1]/a_39_7# mux4_8_10space_0/mux4_dp_1x_0[1]/a_47_7# 2 6 109 121
n inv_1x_8_1/inv_1x_6/y mux4_8_10space_0/mux4_dp_1x_0[1]/a_47_7# mux4_8_10space_0/mux4_dp_1x_0[1]/a_55_7# 2 6 117 121
n op4 mux4_8_10space_0/mux4_dp_1x_0[1]/a_55_7# Gnd! 2 6 122 121
n op3 Gnd! mux4_8_10space_0/mux4_dp_1x_0[1]/a_68_7# 2 6 130 121
n b1 mux4_8_10space_0/mux4_dp_1x_0[1]/a_68_7# mux4_8_10space_0/mux4_dp_1x_0[1]/a_47_7# 2 6 135 121
n mux4_8_10space_0/mux4_dp_1x_0[1]/a_39_7# Gnd! adder_8_0/b_1_ 2 7 157 121
p b2 mux4_8_10space_0/mux4_dp_1x_0[2]/a_6_74# mux4_8_10space_0/mux4_dp_1x_0[2]/a_13_74# 2 9 75 298
p op6 mux4_8_10space_0/mux4_dp_1x_0[2]/a_13_74# Vdd! 2 9 80 298
p op5 Vdd! mux4_8_10space_0/mux4_dp_1x_0[2]/a_26_74# 2 9 88 298
p inv_1x_8_1/inv_1x_5/y mux4_8_10space_0/mux4_dp_1x_0[2]/a_26_74# mux4_8_10space_0/mux4_dp_1x_0[2]/a_6_74# 2 9 93 298
p a2 mux4_8_10space_0/mux4_dp_1x_0[2]/a_6_74# mux4_8_10space_0/mux4_dp_1x_0[2]/a_39_7# 2 9 101 298
p inv_1x_8_0/inv_1x_5/y mux4_8_10space_0/mux4_dp_1x_0[2]/a_39_7# mux4_8_10space_0/mux4_dp_1x_0[2]/a_47_74# 2 9 109 298
p b2 mux4_8_10space_0/mux4_dp_1x_0[2]/a_47_74# mux4_8_10space_0/mux4_dp_1x_0[2]/a_55_74# 2 9 117 298
p op4 mux4_8_10space_0/mux4_dp_1x_0[2]/a_55_74# Vdd! 2 9 122 298
p op3 Vdd! mux4_8_10space_0/mux4_dp_1x_0[2]/a_68_74# 2 9 130 298
p inv_1x_8_1/inv_1x_5/y mux4_8_10space_0/mux4_dp_1x_0[2]/a_68_74# mux4_8_10space_0/mux4_dp_1x_0[2]/a_47_74# 2 9 135 298
p mux4_8_10space_0/mux4_dp_1x_0[2]/a_39_7# Vdd! adder_8_0/b_2_ 2 10 157 297
n inv_1x_8_1/inv_1x_5/y mux4_8_10space_0/mux4_dp_1x_0[2]/a_6_7# mux4_8_10space_0/mux4_dp_1x_0[2]/a_13_7# 2 6 75 231
n op6 mux4_8_10space_0/mux4_dp_1x_0[2]/a_13_7# Gnd! 2 6 80 231
n op5 Gnd! mux4_8_10space_0/mux4_dp_1x_0[2]/a_26_7# 2 6 88 231
n b2 mux4_8_10space_0/mux4_dp_1x_0[2]/a_26_7# mux4_8_10space_0/mux4_dp_1x_0[2]/a_6_7# 2 6 93 231
n inv_1x_8_0/inv_1x_5/y mux4_8_10space_0/mux4_dp_1x_0[2]/a_6_7# mux4_8_10space_0/mux4_dp_1x_0[2]/a_39_7# 2 6 101 231
n a2 mux4_8_10space_0/mux4_dp_1x_0[2]/a_39_7# mux4_8_10space_0/mux4_dp_1x_0[2]/a_47_7# 2 6 109 231
n inv_1x_8_1/inv_1x_5/y mux4_8_10space_0/mux4_dp_1x_0[2]/a_47_7# mux4_8_10space_0/mux4_dp_1x_0[2]/a_55_7# 2 6 117 231
n op4 mux4_8_10space_0/mux4_dp_1x_0[2]/a_55_7# Gnd! 2 6 122 231
n op3 Gnd! mux4_8_10space_0/mux4_dp_1x_0[2]/a_68_7# 2 6 130 231
n b2 mux4_8_10space_0/mux4_dp_1x_0[2]/a_68_7# mux4_8_10space_0/mux4_dp_1x_0[2]/a_47_7# 2 6 135 231
n mux4_8_10space_0/mux4_dp_1x_0[2]/a_39_7# Gnd! adder_8_0/b_2_ 2 7 157 231
p b3 mux4_8_10space_0/mux4_dp_1x_0[3]/a_6_74# mux4_8_10space_0/mux4_dp_1x_0[3]/a_13_74# 2 9 75 408
p op6 mux4_8_10space_0/mux4_dp_1x_0[3]/a_13_74# Vdd! 2 9 80 408
p op5 Vdd! mux4_8_10space_0/mux4_dp_1x_0[3]/a_26_74# 2 9 88 408
p inv_1x_8_1/inv_1x_4/y mux4_8_10space_0/mux4_dp_1x_0[3]/a_26_74# mux4_8_10space_0/mux4_dp_1x_0[3]/a_6_74# 2 9 93 408
p a3 mux4_8_10space_0/mux4_dp_1x_0[3]/a_6_74# mux4_8_10space_0/mux4_dp_1x_0[3]/a_39_7# 2 9 101 408
p inv_1x_8_0/inv_1x_4/y mux4_8_10space_0/mux4_dp_1x_0[3]/a_39_7# mux4_8_10space_0/mux4_dp_1x_0[3]/a_47_74# 2 9 109 408
p b3 mux4_8_10space_0/mux4_dp_1x_0[3]/a_47_74# mux4_8_10space_0/mux4_dp_1x_0[3]/a_55_74# 2 9 117 408
p op4 mux4_8_10space_0/mux4_dp_1x_0[3]/a_55_74# Vdd! 2 9 122 408
p op3 Vdd! mux4_8_10space_0/mux4_dp_1x_0[3]/a_68_74# 2 9 130 408
p inv_1x_8_1/inv_1x_4/y mux4_8_10space_0/mux4_dp_1x_0[3]/a_68_74# mux4_8_10space_0/mux4_dp_1x_0[3]/a_47_74# 2 9 135 408
p mux4_8_10space_0/mux4_dp_1x_0[3]/a_39_7# Vdd! adder_8_0/b_3_ 2 10 157 407
n inv_1x_8_1/inv_1x_4/y mux4_8_10space_0/mux4_dp_1x_0[3]/a_6_7# mux4_8_10space_0/mux4_dp_1x_0[3]/a_13_7# 2 6 75 341
n op6 mux4_8_10space_0/mux4_dp_1x_0[3]/a_13_7# Gnd! 2 6 80 341
n op5 Gnd! mux4_8_10space_0/mux4_dp_1x_0[3]/a_26_7# 2 6 88 341
n b3 mux4_8_10space_0/mux4_dp_1x_0[3]/a_26_7# mux4_8_10space_0/mux4_dp_1x_0[3]/a_6_7# 2 6 93 341
n inv_1x_8_0/inv_1x_4/y mux4_8_10space_0/mux4_dp_1x_0[3]/a_6_7# mux4_8_10space_0/mux4_dp_1x_0[3]/a_39_7# 2 6 101 341
n a3 mux4_8_10space_0/mux4_dp_1x_0[3]/a_39_7# mux4_8_10space_0/mux4_dp_1x_0[3]/a_47_7# 2 6 109 341
n inv_1x_8_1/inv_1x_4/y mux4_8_10space_0/mux4_dp_1x_0[3]/a_47_7# mux4_8_10space_0/mux4_dp_1x_0[3]/a_55_7# 2 6 117 341
n op4 mux4_8_10space_0/mux4_dp_1x_0[3]/a_55_7# Gnd! 2 6 122 341
n op3 Gnd! mux4_8_10space_0/mux4_dp_1x_0[3]/a_68_7# 2 6 130 341
n b3 mux4_8_10space_0/mux4_dp_1x_0[3]/a_68_7# mux4_8_10space_0/mux4_dp_1x_0[3]/a_47_7# 2 6 135 341
n mux4_8_10space_0/mux4_dp_1x_0[3]/a_39_7# Gnd! adder_8_0/b_3_ 2 7 157 341
p b4 mux4_8_10space_0/mux4_dp_1x_0[4]/a_6_74# mux4_8_10space_0/mux4_dp_1x_0[4]/a_13_74# 2 9 75 518
p op6 mux4_8_10space_0/mux4_dp_1x_0[4]/a_13_74# Vdd! 2 9 80 518
p op5 Vdd! mux4_8_10space_0/mux4_dp_1x_0[4]/a_26_74# 2 9 88 518
p inv_1x_8_1/inv_1x_3/y mux4_8_10space_0/mux4_dp_1x_0[4]/a_26_74# mux4_8_10space_0/mux4_dp_1x_0[4]/a_6_74# 2 9 93 518
p a4 mux4_8_10space_0/mux4_dp_1x_0[4]/a_6_74# mux4_8_10space_0/mux4_dp_1x_0[4]/a_39_7# 2 9 101 518
p inv_1x_8_0/inv_1x_3/y mux4_8_10space_0/mux4_dp_1x_0[4]/a_39_7# mux4_8_10space_0/mux4_dp_1x_0[4]/a_47_74# 2 9 109 518
p b4 mux4_8_10space_0/mux4_dp_1x_0[4]/a_47_74# mux4_8_10space_0/mux4_dp_1x_0[4]/a_55_74# 2 9 117 518
p op4 mux4_8_10space_0/mux4_dp_1x_0[4]/a_55_74# Vdd! 2 9 122 518
p op3 Vdd! mux4_8_10space_0/mux4_dp_1x_0[4]/a_68_74# 2 9 130 518
p inv_1x_8_1/inv_1x_3/y mux4_8_10space_0/mux4_dp_1x_0[4]/a_68_74# mux4_8_10space_0/mux4_dp_1x_0[4]/a_47_74# 2 9 135 518
p mux4_8_10space_0/mux4_dp_1x_0[4]/a_39_7# Vdd! adder_8_0/b_4_ 2 10 157 517
n inv_1x_8_1/inv_1x_3/y mux4_8_10space_0/mux4_dp_1x_0[4]/a_6_7# mux4_8_10space_0/mux4_dp_1x_0[4]/a_13_7# 2 6 75 451
n op6 mux4_8_10space_0/mux4_dp_1x_0[4]/a_13_7# Gnd! 2 6 80 451
n op5 Gnd! mux4_8_10space_0/mux4_dp_1x_0[4]/a_26_7# 2 6 88 451
n b4 mux4_8_10space_0/mux4_dp_1x_0[4]/a_26_7# mux4_8_10space_0/mux4_dp_1x_0[4]/a_6_7# 2 6 93 451
n inv_1x_8_0/inv_1x_3/y mux4_8_10space_0/mux4_dp_1x_0[4]/a_6_7# mux4_8_10space_0/mux4_dp_1x_0[4]/a_39_7# 2 6 101 451
n a4 mux4_8_10space_0/mux4_dp_1x_0[4]/a_39_7# mux4_8_10space_0/mux4_dp_1x_0[4]/a_47_7# 2 6 109 451
n inv_1x_8_1/inv_1x_3/y mux4_8_10space_0/mux4_dp_1x_0[4]/a_47_7# mux4_8_10space_0/mux4_dp_1x_0[4]/a_55_7# 2 6 117 451
n op4 mux4_8_10space_0/mux4_dp_1x_0[4]/a_55_7# Gnd! 2 6 122 451
n op3 Gnd! mux4_8_10space_0/mux4_dp_1x_0[4]/a_68_7# 2 6 130 451
n b4 mux4_8_10space_0/mux4_dp_1x_0[4]/a_68_7# mux4_8_10space_0/mux4_dp_1x_0[4]/a_47_7# 2 6 135 451
n mux4_8_10space_0/mux4_dp_1x_0[4]/a_39_7# Gnd! adder_8_0/b_4_ 2 7 157 451
p b5 mux4_8_10space_0/mux4_dp_1x_0[5]/a_6_74# mux4_8_10space_0/mux4_dp_1x_0[5]/a_13_74# 2 9 75 628
p op6 mux4_8_10space_0/mux4_dp_1x_0[5]/a_13_74# Vdd! 2 9 80 628
p op5 Vdd! mux4_8_10space_0/mux4_dp_1x_0[5]/a_26_74# 2 9 88 628
p inv_1x_8_1/inv_1x_2/y mux4_8_10space_0/mux4_dp_1x_0[5]/a_26_74# mux4_8_10space_0/mux4_dp_1x_0[5]/a_6_74# 2 9 93 628
p a5 mux4_8_10space_0/mux4_dp_1x_0[5]/a_6_74# mux4_8_10space_0/mux4_dp_1x_0[5]/a_39_7# 2 9 101 628
p inv_1x_8_0/inv_1x_2/y mux4_8_10space_0/mux4_dp_1x_0[5]/a_39_7# mux4_8_10space_0/mux4_dp_1x_0[5]/a_47_74# 2 9 109 628
p b5 mux4_8_10space_0/mux4_dp_1x_0[5]/a_47_74# mux4_8_10space_0/mux4_dp_1x_0[5]/a_55_74# 2 9 117 628
p op4 mux4_8_10space_0/mux4_dp_1x_0[5]/a_55_74# Vdd! 2 9 122 628
p op3 Vdd! mux4_8_10space_0/mux4_dp_1x_0[5]/a_68_74# 2 9 130 628
p inv_1x_8_1/inv_1x_2/y mux4_8_10space_0/mux4_dp_1x_0[5]/a_68_74# mux4_8_10space_0/mux4_dp_1x_0[5]/a_47_74# 2 9 135 628
p mux4_8_10space_0/mux4_dp_1x_0[5]/a_39_7# Vdd! adder_8_0/b_5_ 2 10 157 627
n inv_1x_8_1/inv_1x_2/y mux4_8_10space_0/mux4_dp_1x_0[5]/a_6_7# mux4_8_10space_0/mux4_dp_1x_0[5]/a_13_7# 2 6 75 561
n op6 mux4_8_10space_0/mux4_dp_1x_0[5]/a_13_7# Gnd! 2 6 80 561
n op5 Gnd! mux4_8_10space_0/mux4_dp_1x_0[5]/a_26_7# 2 6 88 561
n b5 mux4_8_10space_0/mux4_dp_1x_0[5]/a_26_7# mux4_8_10space_0/mux4_dp_1x_0[5]/a_6_7# 2 6 93 561
n inv_1x_8_0/inv_1x_2/y mux4_8_10space_0/mux4_dp_1x_0[5]/a_6_7# mux4_8_10space_0/mux4_dp_1x_0[5]/a_39_7# 2 6 101 561
n a5 mux4_8_10space_0/mux4_dp_1x_0[5]/a_39_7# mux4_8_10space_0/mux4_dp_1x_0[5]/a_47_7# 2 6 109 561
n inv_1x_8_1/inv_1x_2/y mux4_8_10space_0/mux4_dp_1x_0[5]/a_47_7# mux4_8_10space_0/mux4_dp_1x_0[5]/a_55_7# 2 6 117 561
n op4 mux4_8_10space_0/mux4_dp_1x_0[5]/a_55_7# Gnd! 2 6 122 561
n op3 Gnd! mux4_8_10space_0/mux4_dp_1x_0[5]/a_68_7# 2 6 130 561
n b5 mux4_8_10space_0/mux4_dp_1x_0[5]/a_68_7# mux4_8_10space_0/mux4_dp_1x_0[5]/a_47_7# 2 6 135 561
n mux4_8_10space_0/mux4_dp_1x_0[5]/a_39_7# Gnd! adder_8_0/b_5_ 2 7 157 561
p b6 mux4_8_10space_0/mux4_dp_1x_0[6]/a_6_74# mux4_8_10space_0/mux4_dp_1x_0[6]/a_13_74# 2 9 75 738
p op6 mux4_8_10space_0/mux4_dp_1x_0[6]/a_13_74# Vdd! 2 9 80 738
p op5 Vdd! mux4_8_10space_0/mux4_dp_1x_0[6]/a_26_74# 2 9 88 738
p inv_1x_8_1/inv_1x_1/y mux4_8_10space_0/mux4_dp_1x_0[6]/a_26_74# mux4_8_10space_0/mux4_dp_1x_0[6]/a_6_74# 2 9 93 738
p a6 mux4_8_10space_0/mux4_dp_1x_0[6]/a_6_74# mux4_8_10space_0/mux4_dp_1x_0[6]/a_39_7# 2 9 101 738
p inv_1x_8_0/inv_1x_1/y mux4_8_10space_0/mux4_dp_1x_0[6]/a_39_7# mux4_8_10space_0/mux4_dp_1x_0[6]/a_47_74# 2 9 109 738
p b6 mux4_8_10space_0/mux4_dp_1x_0[6]/a_47_74# mux4_8_10space_0/mux4_dp_1x_0[6]/a_55_74# 2 9 117 738
p op4 mux4_8_10space_0/mux4_dp_1x_0[6]/a_55_74# Vdd! 2 9 122 738
p op3 Vdd! mux4_8_10space_0/mux4_dp_1x_0[6]/a_68_74# 2 9 130 738
p inv_1x_8_1/inv_1x_1/y mux4_8_10space_0/mux4_dp_1x_0[6]/a_68_74# mux4_8_10space_0/mux4_dp_1x_0[6]/a_47_74# 2 9 135 738
p mux4_8_10space_0/mux4_dp_1x_0[6]/a_39_7# Vdd! adder_8_0/b_6_ 2 10 157 737
n inv_1x_8_1/inv_1x_1/y mux4_8_10space_0/mux4_dp_1x_0[6]/a_6_7# mux4_8_10space_0/mux4_dp_1x_0[6]/a_13_7# 2 6 75 671
n op6 mux4_8_10space_0/mux4_dp_1x_0[6]/a_13_7# Gnd! 2 6 80 671
n op5 Gnd! mux4_8_10space_0/mux4_dp_1x_0[6]/a_26_7# 2 6 88 671
n b6 mux4_8_10space_0/mux4_dp_1x_0[6]/a_26_7# mux4_8_10space_0/mux4_dp_1x_0[6]/a_6_7# 2 6 93 671
n inv_1x_8_0/inv_1x_1/y mux4_8_10space_0/mux4_dp_1x_0[6]/a_6_7# mux4_8_10space_0/mux4_dp_1x_0[6]/a_39_7# 2 6 101 671
n a6 mux4_8_10space_0/mux4_dp_1x_0[6]/a_39_7# mux4_8_10space_0/mux4_dp_1x_0[6]/a_47_7# 2 6 109 671
n inv_1x_8_1/inv_1x_1/y mux4_8_10space_0/mux4_dp_1x_0[6]/a_47_7# mux4_8_10space_0/mux4_dp_1x_0[6]/a_55_7# 2 6 117 671
n op4 mux4_8_10space_0/mux4_dp_1x_0[6]/a_55_7# Gnd! 2 6 122 671
n op3 Gnd! mux4_8_10space_0/mux4_dp_1x_0[6]/a_68_7# 2 6 130 671
n b6 mux4_8_10space_0/mux4_dp_1x_0[6]/a_68_7# mux4_8_10space_0/mux4_dp_1x_0[6]/a_47_7# 2 6 135 671
n mux4_8_10space_0/mux4_dp_1x_0[6]/a_39_7# Gnd! adder_8_0/b_6_ 2 7 157 671
p b7 mux4_8_10space_0/mux4_dp_1x_0[7]/a_6_74# mux4_8_10space_0/mux4_dp_1x_0[7]/a_13_74# 2 9 75 848
p op6 mux4_8_10space_0/mux4_dp_1x_0[7]/a_13_74# Vdd! 2 9 80 848
p op5 Vdd! mux4_8_10space_0/mux4_dp_1x_0[7]/a_26_74# 2 9 88 848
p inv_1x_8_1/inv_1x_0/y mux4_8_10space_0/mux4_dp_1x_0[7]/a_26_74# mux4_8_10space_0/mux4_dp_1x_0[7]/a_6_74# 2 9 93 848
p a7 mux4_8_10space_0/mux4_dp_1x_0[7]/a_6_74# mux4_8_10space_0/mux4_dp_1x_0[7]/a_39_7# 2 9 101 848
p inv_1x_8_0/inv_1x_0/y mux4_8_10space_0/mux4_dp_1x_0[7]/a_39_7# mux4_8_10space_0/mux4_dp_1x_0[7]/a_47_74# 2 9 109 848
p b7 mux4_8_10space_0/mux4_dp_1x_0[7]/a_47_74# mux4_8_10space_0/mux4_dp_1x_0[7]/a_55_74# 2 9 117 848
p op4 mux4_8_10space_0/mux4_dp_1x_0[7]/a_55_74# Vdd! 2 9 122 848
p op3 Vdd! mux4_8_10space_0/mux4_dp_1x_0[7]/a_68_74# 2 9 130 848
p inv_1x_8_1/inv_1x_0/y mux4_8_10space_0/mux4_dp_1x_0[7]/a_68_74# mux4_8_10space_0/mux4_dp_1x_0[7]/a_47_74# 2 9 135 848
p mux4_8_10space_0/mux4_dp_1x_0[7]/a_39_7# Vdd! adder_8_0/b_7_ 2 10 157 847
n inv_1x_8_1/inv_1x_0/y mux4_8_10space_0/mux4_dp_1x_0[7]/a_6_7# mux4_8_10space_0/mux4_dp_1x_0[7]/a_13_7# 2 6 75 781
n op6 mux4_8_10space_0/mux4_dp_1x_0[7]/a_13_7# Gnd! 2 6 80 781
n op5 Gnd! mux4_8_10space_0/mux4_dp_1x_0[7]/a_26_7# 2 6 88 781
n b7 mux4_8_10space_0/mux4_dp_1x_0[7]/a_26_7# mux4_8_10space_0/mux4_dp_1x_0[7]/a_6_7# 2 6 93 781
n inv_1x_8_0/inv_1x_0/y mux4_8_10space_0/mux4_dp_1x_0[7]/a_6_7# mux4_8_10space_0/mux4_dp_1x_0[7]/a_39_7# 2 6 101 781
n a7 mux4_8_10space_0/mux4_dp_1x_0[7]/a_39_7# mux4_8_10space_0/mux4_dp_1x_0[7]/a_47_7# 2 6 109 781
n inv_1x_8_1/inv_1x_0/y mux4_8_10space_0/mux4_dp_1x_0[7]/a_47_7# mux4_8_10space_0/mux4_dp_1x_0[7]/a_55_7# 2 6 117 781
n op4 mux4_8_10space_0/mux4_dp_1x_0[7]/a_55_7# Gnd! 2 6 122 781
n op3 Gnd! mux4_8_10space_0/mux4_dp_1x_0[7]/a_68_7# 2 6 130 781
n b7 mux4_8_10space_0/mux4_dp_1x_0[7]/a_68_7# mux4_8_10space_0/mux4_dp_1x_0[7]/a_47_7# 2 6 135 781
n mux4_8_10space_0/mux4_dp_1x_0[7]/a_39_7# Gnd! adder_8_0/b_7_ 2 7 157 781
p b0 Vdd! inv_1x_8_1/inv_1x_7/y 2 10 53 77
n b0 Gnd! inv_1x_8_1/inv_1x_7/y 2 7 53 11
p b1 Vdd! inv_1x_8_1/inv_1x_6/y 2 10 53 187
n b1 Gnd! inv_1x_8_1/inv_1x_6/y 2 7 53 121
p b2 Vdd! inv_1x_8_1/inv_1x_5/y 2 10 53 297
n b2 Gnd! inv_1x_8_1/inv_1x_5/y 2 7 53 231
p b3 Vdd! inv_1x_8_1/inv_1x_4/y 2 10 53 407
n b3 Gnd! inv_1x_8_1/inv_1x_4/y 2 7 53 341
p b4 Vdd! inv_1x_8_1/inv_1x_3/y 2 10 53 517
n b4 Gnd! inv_1x_8_1/inv_1x_3/y 2 7 53 451
p b5 Vdd! inv_1x_8_1/inv_1x_2/y 2 10 53 627
n b5 Gnd! inv_1x_8_1/inv_1x_2/y 2 7 53 561
p b6 Vdd! inv_1x_8_1/inv_1x_1/y 2 10 53 737
n b6 Gnd! inv_1x_8_1/inv_1x_1/y 2 7 53 671
p b7 Vdd! inv_1x_8_1/inv_1x_0/y 2 10 53 847
n b7 Gnd! inv_1x_8_1/inv_1x_0/y 2 7 53 781
p a0 Vdd! inv_1x_8_0/inv_1x_7/y 2 10 37 77
n a0 Gnd! inv_1x_8_0/inv_1x_7/y 2 7 37 11
p a1 Vdd! inv_1x_8_0/inv_1x_6/y 2 10 37 187
n a1 Gnd! inv_1x_8_0/inv_1x_6/y 2 7 37 121
p a2 Vdd! inv_1x_8_0/inv_1x_5/y 2 10 37 297
n a2 Gnd! inv_1x_8_0/inv_1x_5/y 2 7 37 231
p a3 Vdd! inv_1x_8_0/inv_1x_4/y 2 10 37 407
n a3 Gnd! inv_1x_8_0/inv_1x_4/y 2 7 37 341
p a4 Vdd! inv_1x_8_0/inv_1x_3/y 2 10 37 517
n a4 Gnd! inv_1x_8_0/inv_1x_3/y 2 7 37 451
p a5 Vdd! inv_1x_8_0/inv_1x_2/y 2 10 37 627
n a5 Gnd! inv_1x_8_0/inv_1x_2/y 2 7 37 561
p a6 Vdd! inv_1x_8_0/inv_1x_1/y 2 10 37 737
n a6 Gnd! inv_1x_8_0/inv_1x_1/y 2 7 37 671
p a7 Vdd! inv_1x_8_0/inv_1x_0/y 2 10 37 847
n a7 Gnd! inv_1x_8_0/inv_1x_0/y 2 7 37 781
p result0 Vdd! yzdetect_8_0/nor2_1x_4/a_7_67# 2 16 5 71
p result1 yzdetect_8_0/nor2_1x_4/a_7_67# yzdetect_8_0/nor2_1x_4/y 2 16 10 71
n result0 Gnd! yzdetect_8_0/nor2_1x_4/y 2 8 5 11
n result1 yzdetect_8_0/nor2_1x_4/y Gnd! 2 8 13 11
p yzdetect_8_0/nor2_1x_4/y Vdd! yzdetect_8_0/nor2_1x_2/b 2 12 5 185
p yzdetect_8_0/nor2_1x_3/y yzdetect_8_0/nor2_1x_2/b Vdd! 2 12 13 185
n yzdetect_8_0/nor2_1x_4/y Gnd! yzdetect_8_0/nand2_1x_1/a_7_7# 2 12 5 121
n yzdetect_8_0/nor2_1x_3/y yzdetect_8_0/nand2_1x_1/a_7_7# yzdetect_8_0/nor2_1x_2/b 2 12 10 121
p result2 Vdd! yzdetect_8_0/nor2_1x_3/a_7_67# 2 16 5 291
p result3 yzdetect_8_0/nor2_1x_3/a_7_67# yzdetect_8_0/nor2_1x_3/y 2 16 10 291
n result2 Gnd! yzdetect_8_0/nor2_1x_3/y 2 8 5 231
n result3 yzdetect_8_0/nor2_1x_3/y Gnd! 2 8 13 231
p yzdetect_8_0/nor2_1x_2/a Vdd! yzdetect_8_0/nor2_1x_2/a_7_67# 2 16 5 401
p yzdetect_8_0/nor2_1x_2/b yzdetect_8_0/nor2_1x_2/a_7_67# zero 2 16 10 401
n yzdetect_8_0/nor2_1x_2/a Gnd! zero 2 8 5 341
n yzdetect_8_0/nor2_1x_2/b zero Gnd! 2 8 13 341
p result4 Vdd! yzdetect_8_0/nor2_1x_1/a_7_67# 2 16 5 511
p result5 yzdetect_8_0/nor2_1x_1/a_7_67# yzdetect_8_0/nor2_1x_1/y 2 16 10 511
n result4 Gnd! yzdetect_8_0/nor2_1x_1/y 2 8 5 451
n result5 yzdetect_8_0/nor2_1x_1/y Gnd! 2 8 13 451
p yzdetect_8_0/nor2_1x_0/y Vdd! yzdetect_8_0/nor2_1x_2/a 2 12 5 625
p yzdetect_8_0/nor2_1x_1/y yzdetect_8_0/nor2_1x_2/a Vdd! 2 12 13 625
n yzdetect_8_0/nor2_1x_0/y Gnd! yzdetect_8_0/nand2_1x_0/a_7_7# 2 12 5 561
n yzdetect_8_0/nor2_1x_1/y yzdetect_8_0/nand2_1x_0/a_7_7# yzdetect_8_0/nor2_1x_2/a 2 12 10 561
p result6 Vdd! yzdetect_8_0/nor2_1x_0/a_7_67# 2 16 5 731
p result7 yzdetect_8_0/nor2_1x_0/a_7_67# yzdetect_8_0/nor2_1x_0/y 2 16 10 731
n result6 Gnd! yzdetect_8_0/nor2_1x_0/y 2 8 5 671
n result7 yzdetect_8_0/nor2_1x_0/y Gnd! 2 8 13 671
p cout_adder_7 Vdd! inv_1x_0/y 2 10 270 957
n cout_adder_7 Gnd! inv_1x_0/y 2 7 270 891
C Vdd! a4 4.4
C result5 mux3_1x_8_0/mux3_dp_1x_2/a_33_7# 2.1
C Vdd! op5 8.6
C Vdd! alu_ctl_0/OAI21X1_6/C 3.1
C Vdd! adder_8_0/s_4_ 2.6
C Vdd! alu_ctl_0/NAND3X1_0/Y 6.5
C Vdd! adder_8_0/c_7_ 10.4
C Vdd! muxy7 7.1
C Vdd! mux3_1x_8_0/mux3_dp_1x_3/a_0_74# 2.2
C Vdd! adder_8_0/c_6_ 10.4
C Vdd! mux3_1x_8_0/mux3_dp_1x_7/s0b 13.3
C Vdd! alu_ctl_0/NAND3X1_2/Y 5.4
C Vdd! mux3_1x_8_0/mux3_dp_1x_0/a_33_7# 3.1
C Vdd! adder_8_0/b_5_ 7.1
C Vdd! alu_ctl_0/OR2X1_0/a_2_54# 2.1
C Vdd! inv_1x_8_0/inv_1x_6/y 2.7
C Vdd! result1 2.2
C Vdd! op1 2.8
C Vdd! mux3_1x_8_0/mux3_dp_1x_5/a_0_74# 2.2
C Vdd! alu_ctl_0/OAI21X1_2/B 2.0
C Vdd! inv_1x_8_0/inv_1x_0/y 2.7
C result2 mux3_1x_8_0/mux3_dp_1x_5/a_33_7# 2.1
C Vdd! adder_8_0/b_7_ 7.1
C Vdd! op2 7.2
C Vdd! mux3_1x_8_0/mux3_dp_1x_0/a_0_74# 2.2
C Vdd! yzdetect_8_0/nor2_1x_4/y 2.5
C Vdd! alu_ctl_0/INVX2_2/Y 3.5
C Vdd! yzdetect_8_0/nor2_1x_3/y 3.3
C Vdd! inv_1x_8_0/inv_1x_3/y 2.7
C Vdd! b7 6.0
C Vdd! mux3_1x_8_0/mux3_dp_1x_2/a_33_7# 3.1
C Vdd! adder_8_0/b_4_ 7.1
C Vdd! alu_op_1 5.2
C Vdd! mux3_1x_8_0/mux3_dp_1x_1/a_33_7# 3.1
C Vdd! funct_1 7.7
C Vdd! mux3_1x_8_0/mux3_dp_1x_4/a_0_74# 2.2
C Vdd! inv_1x_8_0/inv_1x_5/y 2.7
C a3 Vdd! 4.4
C Vdd! alu_ctl_0/INVX2_3/A 3.5
C Vdd! inv_1x_8_1/inv_1x_6/y 7.0
C Vdd! mux3_1x_8_0/mux3_dp_1x_5/a_33_7# 3.1
C Vdd! adder_8_0/b_6_ 7.1
C Vdd! inv_1x_8_0/inv_1x_1/y 2.7
C Vdd! alu_ctl_0/INVX2_3/Y 3.2
C Vdd! mux3_1x_8_0/mux3_dp_1x_7/a_0_74# 2.2
C Vdd! alu_ctl_0/INVX2_6/Y 2.6
C inv_1x_8_0/inv_1x_2/y Vdd! 2.7
C Vdd! adder_8_0/s_5_ 2.6
C Vdd! mux3_1x_8_0/mux3_dp_1x_4/a_33_7# 3.1
C Vdd! funct_0 5.6
C Vdd! alu_ctl_0/NOR2X1_0/Y 2.8
C Vdd! less 10.9
C yzdetect_8_0/nor2_1x_1/y Vdd! 3.2
C Vdd! op3 8.8
C Vdd! mux3_1x_8_0/mux3_dp_1x_2/a_0_74# 2.2
C Vdd! mux3_1x_8_0/mux3_dp_1x_7/s1b 13.3
C Vdd! alu_ctl_0/AND2X2_0/Y 3.0
C Vdd! b2 5.9
C Vdd! mux3_1x_8_0/mux3_dp_1x_3/a_33_7# 3.1
C Vdd! alu_ctl_0/INVX2_5/Y 3.0
C Vdd! alu_ctl_0/NOR2X1_0/A 3.5
C Vdd! result4 2.5
C Vdd! adder_8_0/s_0_ 2.6
C a6 Vdd! 4.4
C Vdd! inv_1x_8_0/inv_1x_4/y 2.7
C yzdetect_8_0/nor2_1x_0/y Vdd! 2.7
C Vdd! a5 4.4
C Vdd! adder_8_0/c_3_ 10.4
C Vdd! adder_8_0/b_1_ 7.1
C Vdd! yzdetect_8_0/nor2_1x_2/a 3.5
C result0 mux3_1x_8_0/mux3_dp_1x_7/a_33_7# 2.1
C inv_1x_8_1/inv_1x_1/y Vdd! 7.0
C Vdd! op6 8.5
C Vdd! adder_8_0/b_3_ 7.1
C Vdd! alu_ctl_0/OR2X1_0/Y 2.8
C Vdd! result6 2.5
C Vdd! b5 5.9
C Vdd! alu_ctl_0/OAI21X1_7/A 2.4
C Vdd! op0 4.1
C Vdd! result3 2.2
C Vdd! b6 5.9
C Vdd! funct_3 3.1
C Vdd! mux3_1x_8_0/mux3_dp_1x_7/s1 14.0
C Vdd! alu_ctl_0/OAI21X1_7/B 3.2
C Vdd! alu_ctl_0/NOR2X1_2/Y 4.0
C Vdd! inv_1x_8_1/inv_1x_5/y 7.0
C Vdd! adder_8_0/c_1_ 10.4
C Vdd! adder_8_0/s_7_ 2.6
C Vdd! adder_8_0/s_1_ 2.6
C Vdd! inv_1x_8_1/inv_1x_7/y 7.0
C Vdd! alu_ctl_0/OAI21X1_2/C 5.7
C Vdd! inv_1x_0/y 5.0
C Vdd! op4 15.4
C Vdd! inv_1x_8_1/inv_1x_0/y 7.0
C Vdd! adder_8_0/c_4_ 10.4
C adder_8_0/s_2_ Vdd! 2.6
C Vdd! mux3_1x_8_0/mux3_dp_1x_7/a_33_7# 3.1
C Vdd! a7 4.4
C Vdd! adder_8_0/s_6_ 2.6
C Vdd! funct_2 3.7
C Vdd! inv_1x_8_1/inv_1x_4/y 7.0
C Vdd! adder_8_0/c_5_ 10.4
C a2 Vdd! 4.4
C Vdd! mux3_1x_8_0/mux3_dp_1x_6/a_33_7# 3.1
C Vdd! alu_ctl_0/INVX2_1/A 6.0
C result6 mux3_1x_8_0/mux3_dp_1x_1/a_33_7# 2.1
C Vdd! adder_8_0/s_3_ 2.6
C Vdd! b0 5.9
C result7 mux3_1x_8_0/mux3_dp_1x_0/a_33_7# 2.1
C Vdd! a0 4.4
C Vdd! result7 2.2
C result1 mux3_1x_8_0/mux3_dp_1x_6/a_33_7# 2.1
C Vdd! b4 5.9
C inv_1x_8_0/inv_1x_7/y Vdd! 2.7
C result4 mux3_1x_8_0/mux3_dp_1x_3/a_33_7# 2.1
C Vdd! alu_ctl_0/NAND2X1_5/B 2.4
C Vdd! result5 2.7
C Vdd! alu_op_0 4.2
C yzdetect_8_0/nor2_1x_2/b Vdd! 3.2
C Vdd! adder_8_0/c_2_ 10.4
C Vdd! mux3_1x_8_0/mux3_dp_1x_7/s0 11.5
C Vdd! inv_1x_8_1/inv_1x_2/y 7.0
C Vdd! b3 5.9
C Vdd! adder_8_0/b_2_ 7.1
C Vdd! alu_ctl_0/INVX2_0/Y 5.2
C mux3_1x_8_0/mux3_dp_1x_4/a_33_7# result3 2.1
C Vdd! mux3_1x_8_0/mux3_dp_1x_6/a_0_74# 2.2
C Vdd! result0 2.5
C Vdd! result2 2.5
C Vdd! a1 4.4
C Vdd! alu_ctl_0/INVX2_4/Y 2.9
C Vdd! inv_1x_8_1/inv_1x_3/y 7.0
C mux3_1x_8_0/mux3_dp_1x_7/s1 mux3_1x_8_0/mux3_dp_1x_7/s1b 2.8
C Vdd! b1 5.9
C Vdd! mux3_1x_8_0/mux3_dp_1x_1/a_0_74# 2.2
C Vdd! cout_adder_7 7.0
C inv_1x_0/y GND 7.4
R inv_1x_0/y 1590
C cout_adder_7 GND 7.8
R cout_adder_7 1356
C yzdetect_8_0/nor2_1x_0/y GND 6.7
R yzdetect_8_0/nor2_1x_0/y 1332
R yzdetect_8_0/nor2_1x_0/a_7_67# 561
R yzdetect_8_0/nand2_1x_0/a_7_7# 329
C yzdetect_8_0/nor2_1x_2/a GND 7.3
R yzdetect_8_0/nor2_1x_2/a 1294
C yzdetect_8_0/nor2_1x_1/y GND 7.0
R yzdetect_8_0/nor2_1x_1/y 1365
R yzdetect_8_0/nor2_1x_1/a_7_67# 561
R zero 448
R yzdetect_8_0/nor2_1x_2/a_7_67# 561
C yzdetect_8_0/nor2_1x_2/b GND 7.3
R yzdetect_8_0/nor2_1x_2/b 1326
C yzdetect_8_0/nor2_1x_3/y GND 5.7
R yzdetect_8_0/nor2_1x_3/y 1364
R yzdetect_8_0/nor2_1x_3/a_7_67# 561
R yzdetect_8_0/nand2_1x_1/a_7_7# 329
C yzdetect_8_0/nor2_1x_4/y GND 7.2
R yzdetect_8_0/nor2_1x_4/y 1332
R yzdetect_8_0/nor2_1x_4/a_7_67# 561
C inv_1x_8_0/inv_1x_0/y GND 5.8
R inv_1x_8_0/inv_1x_0/y 1335
R mux4_8_10space_0/mux4_dp_1x_0[7]/a_68_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[7]/a_55_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[7]/a_47_7# 481
R mux4_8_10space_0/mux4_dp_1x_0[7]/a_26_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[7]/a_13_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[7]/a_6_7# 481
R mux4_8_10space_0/mux4_dp_1x_0[7]/a_68_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[7]/a_55_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[7]/a_47_74# 668
R mux4_8_10space_0/mux4_dp_1x_0[7]/a_26_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[7]/a_13_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[7]/a_6_74# 668
C mux4_8_10space_0/mux4_dp_1x_0[7]/a_39_7# GND 3.8
R mux4_8_10space_0/mux4_dp_1x_0[7]/a_39_7# 1123
C op3 GND 44.2
R op3 9028
C op4 GND 47.8
R op4 9068
C a7 GND 11.2
R a7 5505
C inv_1x_8_1/inv_1x_0/y GND 3.3
R inv_1x_8_1/inv_1x_0/y 2524
C op5 GND 42.9
R op5 8846
C op6 GND 43.5
R op6 8489
C b7 GND 6.2
R b7 3063
R mux4_8_10space_0/mux4_dp_1x_0[6]/a_68_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[6]/a_55_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[6]/a_47_7# 481
R mux4_8_10space_0/mux4_dp_1x_0[6]/a_26_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[6]/a_13_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[6]/a_6_7# 481
R mux4_8_10space_0/mux4_dp_1x_0[6]/a_68_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[6]/a_55_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[6]/a_47_74# 668
R mux4_8_10space_0/mux4_dp_1x_0[6]/a_26_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[6]/a_13_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[6]/a_6_74# 668
C mux4_8_10space_0/mux4_dp_1x_0[6]/a_39_7# GND 3.8
R mux4_8_10space_0/mux4_dp_1x_0[6]/a_39_7# 1123
C inv_1x_8_0/inv_1x_1/y GND 5.5
R inv_1x_8_0/inv_1x_1/y 1335
C a6 GND 10.7
R a6 5505
C inv_1x_8_1/inv_1x_1/y GND 3.3
R inv_1x_8_1/inv_1x_1/y 2525
C b6 GND 5.8
R b6 3064
R mux4_8_10space_0/mux4_dp_1x_0[5]/a_68_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[5]/a_55_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[5]/a_47_7# 481
R mux4_8_10space_0/mux4_dp_1x_0[5]/a_26_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[5]/a_13_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[5]/a_6_7# 481
R mux4_8_10space_0/mux4_dp_1x_0[5]/a_68_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[5]/a_55_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[5]/a_47_74# 668
R mux4_8_10space_0/mux4_dp_1x_0[5]/a_26_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[5]/a_13_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[5]/a_6_74# 668
C mux4_8_10space_0/mux4_dp_1x_0[5]/a_39_7# GND 3.8
R mux4_8_10space_0/mux4_dp_1x_0[5]/a_39_7# 1123
C inv_1x_8_0/inv_1x_2/y GND 5.6
R inv_1x_8_0/inv_1x_2/y 1335
C inv_1x_8_1/inv_1x_2/y GND 3.3
R inv_1x_8_1/inv_1x_2/y 2525
C b5 GND 5.8
R b5 3063
R mux4_8_10space_0/mux4_dp_1x_0[4]/a_68_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[4]/a_55_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[4]/a_47_7# 481
R mux4_8_10space_0/mux4_dp_1x_0[4]/a_26_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[4]/a_13_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[4]/a_6_7# 481
R mux4_8_10space_0/mux4_dp_1x_0[4]/a_68_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[4]/a_55_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[4]/a_47_74# 668
R mux4_8_10space_0/mux4_dp_1x_0[4]/a_26_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[4]/a_13_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[4]/a_6_74# 668
C mux4_8_10space_0/mux4_dp_1x_0[4]/a_39_7# GND 3.8
R mux4_8_10space_0/mux4_dp_1x_0[4]/a_39_7# 1123
C inv_1x_8_0/inv_1x_3/y GND 5.5
R inv_1x_8_0/inv_1x_3/y 1335
C inv_1x_8_1/inv_1x_3/y GND 3.3
R inv_1x_8_1/inv_1x_3/y 2524
C b4 GND 4.4
R b4 3063
R mux4_8_10space_0/mux4_dp_1x_0[3]/a_68_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[3]/a_55_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[3]/a_47_7# 481
R mux4_8_10space_0/mux4_dp_1x_0[3]/a_26_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[3]/a_13_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[3]/a_6_7# 481
R mux4_8_10space_0/mux4_dp_1x_0[3]/a_68_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[3]/a_55_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[3]/a_47_74# 668
R mux4_8_10space_0/mux4_dp_1x_0[3]/a_26_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[3]/a_13_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[3]/a_6_74# 668
C mux4_8_10space_0/mux4_dp_1x_0[3]/a_39_7# GND 3.8
R mux4_8_10space_0/mux4_dp_1x_0[3]/a_39_7# 1123
C inv_1x_8_0/inv_1x_4/y GND 5.5
R inv_1x_8_0/inv_1x_4/y 1335
C inv_1x_8_1/inv_1x_4/y GND 3.3
R inv_1x_8_1/inv_1x_4/y 2524
C b3 GND 6.4
R b3 3063
R mux4_8_10space_0/mux4_dp_1x_0[2]/a_68_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[2]/a_55_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[2]/a_47_7# 481
R mux4_8_10space_0/mux4_dp_1x_0[2]/a_26_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[2]/a_13_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[2]/a_6_7# 481
R mux4_8_10space_0/mux4_dp_1x_0[2]/a_68_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[2]/a_55_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[2]/a_47_74# 668
R mux4_8_10space_0/mux4_dp_1x_0[2]/a_26_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[2]/a_13_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[2]/a_6_74# 668
C mux4_8_10space_0/mux4_dp_1x_0[2]/a_39_7# GND 3.8
R mux4_8_10space_0/mux4_dp_1x_0[2]/a_39_7# 1123
C inv_1x_8_0/inv_1x_5/y GND 5.5
R inv_1x_8_0/inv_1x_5/y 1335
C inv_1x_8_1/inv_1x_5/y GND 3.3
R inv_1x_8_1/inv_1x_5/y 2524
C b2 GND 5.8
R b2 3063
R mux4_8_10space_0/mux4_dp_1x_0[1]/a_68_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[1]/a_55_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[1]/a_47_7# 481
R mux4_8_10space_0/mux4_dp_1x_0[1]/a_26_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[1]/a_13_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[1]/a_6_7# 481
R mux4_8_10space_0/mux4_dp_1x_0[1]/a_68_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[1]/a_55_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[1]/a_47_74# 668
R mux4_8_10space_0/mux4_dp_1x_0[1]/a_26_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[1]/a_13_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[1]/a_6_74# 668
C mux4_8_10space_0/mux4_dp_1x_0[1]/a_39_7# GND 3.8
R mux4_8_10space_0/mux4_dp_1x_0[1]/a_39_7# 1123
C inv_1x_8_0/inv_1x_6/y GND 5.5
R inv_1x_8_0/inv_1x_6/y 1335
C inv_1x_8_1/inv_1x_6/y GND 3.3
R inv_1x_8_1/inv_1x_6/y 2524
C b1 GND 5.8
R b1 3063
R mux4_8_10space_0/mux4_dp_1x_0[0]/a_68_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[0]/a_55_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[0]/a_47_7# 481
R mux4_8_10space_0/mux4_dp_1x_0[0]/a_26_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[0]/a_13_7# 164
R mux4_8_10space_0/mux4_dp_1x_0[0]/a_6_7# 481
R mux4_8_10space_0/mux4_dp_1x_0[0]/a_68_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[0]/a_55_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[0]/a_47_74# 668
R mux4_8_10space_0/mux4_dp_1x_0[0]/a_26_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[0]/a_13_74# 316
R mux4_8_10space_0/mux4_dp_1x_0[0]/a_6_74# 668
C mux4_8_10space_0/mux4_dp_1x_0[0]/a_39_7# GND 3.8
R mux4_8_10space_0/mux4_dp_1x_0[0]/a_39_7# 1123
C inv_1x_8_0/inv_1x_7/y GND 5.7
R inv_1x_8_0/inv_1x_7/y 1335
C inv_1x_8_1/inv_1x_7/y GND 3.3
R inv_1x_8_1/inv_1x_7/y 2524
C b0 GND 5.8
R b0 3063
R adder_8_0/fulladder_0/a_85_7# 110
R adder_8_0/fulladder_0/a_77_7# 110
R adder_8_0/fulladder_0/a_45_7# 494
R adder_8_0/fulladder_0/a_29_7# 110
R adder_8_0/fulladder_0/a_n2_7# 504
R adder_8_0/fulladder_0/a_85_65# 281
R adder_8_0/fulladder_0/a_77_65# 281
R adder_8_0/fulladder_0/a_45_65# 838
R adder_8_0/fulladder_0/a_29_65# 281
R adder_8_0/fulladder_0/a_n2_65# 883
C adder_8_0/fulladder_0/a_69_7# GND 2.4
R adder_8_0/fulladder_0/a_69_7# 1250
C adder_8_0/fulladder_0/a_21_7# GND 5.8
R adder_8_0/fulladder_0/a_21_7# 2154
C adder_8_0/c_7_ GND 5.7
R adder_8_0/c_7_ 3139
R adder_8_0/fulladder_1/a_85_7# 110
R adder_8_0/fulladder_1/a_77_7# 110
R adder_8_0/fulladder_1/a_45_7# 494
R adder_8_0/fulladder_1/a_29_7# 110
R adder_8_0/fulladder_1/a_n2_7# 504
R adder_8_0/fulladder_1/a_85_65# 281
R adder_8_0/fulladder_1/a_77_65# 281
R adder_8_0/fulladder_1/a_45_65# 838
R adder_8_0/fulladder_1/a_29_65# 281
R adder_8_0/fulladder_1/a_n2_65# 883
C adder_8_0/fulladder_1/a_69_7# GND 2.4
R adder_8_0/fulladder_1/a_69_7# 1250
C adder_8_0/fulladder_1/a_21_7# GND 5.8
R adder_8_0/fulladder_1/a_21_7# 2154
C adder_8_0/c_6_ GND 5.7
R adder_8_0/c_6_ 3139
R adder_8_0/fulladder_2/a_85_7# 110
R adder_8_0/fulladder_2/a_77_7# 110
R adder_8_0/fulladder_2/a_45_7# 494
R adder_8_0/fulladder_2/a_29_7# 110
R adder_8_0/fulladder_2/a_n2_7# 504
R adder_8_0/fulladder_2/a_85_65# 281
R adder_8_0/fulladder_2/a_77_65# 281
R adder_8_0/fulladder_2/a_45_65# 838
R adder_8_0/fulladder_2/a_29_65# 281
R adder_8_0/fulladder_2/a_n2_65# 883
C adder_8_0/fulladder_2/a_69_7# GND 2.4
R adder_8_0/fulladder_2/a_69_7# 1250
C adder_8_0/fulladder_2/a_21_7# GND 5.8
R adder_8_0/fulladder_2/a_21_7# 2154
C adder_8_0/c_5_ GND 5.7
R adder_8_0/c_5_ 3139
C a5 GND 10.8
R a5 5505
R adder_8_0/fulladder_3/a_85_7# 110
R adder_8_0/fulladder_3/a_77_7# 110
R adder_8_0/fulladder_3/a_45_7# 494
R adder_8_0/fulladder_3/a_29_7# 110
R adder_8_0/fulladder_3/a_n2_7# 504
R adder_8_0/fulladder_3/a_85_65# 281
R adder_8_0/fulladder_3/a_77_65# 281
R adder_8_0/fulladder_3/a_45_65# 838
R adder_8_0/fulladder_3/a_29_65# 281
R adder_8_0/fulladder_3/a_n2_65# 883
C adder_8_0/fulladder_3/a_69_7# GND 2.4
R adder_8_0/fulladder_3/a_69_7# 1250
C adder_8_0/fulladder_3/a_21_7# GND 5.8
R adder_8_0/fulladder_3/a_21_7# 2154
C adder_8_0/c_4_ GND 5.7
R adder_8_0/c_4_ 3138
C a4 GND 10.8
R a4 5505
R adder_8_0/fulladder_4/a_85_7# 110
R adder_8_0/fulladder_4/a_77_7# 110
R adder_8_0/fulladder_4/a_45_7# 494
R adder_8_0/fulladder_4/a_29_7# 110
R adder_8_0/fulladder_4/a_n2_7# 504
R adder_8_0/fulladder_4/a_85_65# 281
R adder_8_0/fulladder_4/a_77_65# 281
R adder_8_0/fulladder_4/a_45_65# 838
R adder_8_0/fulladder_4/a_29_65# 281
R adder_8_0/fulladder_4/a_n2_65# 883
C adder_8_0/fulladder_4/a_69_7# GND 2.4
R adder_8_0/fulladder_4/a_69_7# 1250
C adder_8_0/fulladder_4/a_21_7# GND 5.8
R adder_8_0/fulladder_4/a_21_7# 2154
C adder_8_0/c_3_ GND 5.7
R adder_8_0/c_3_ 3139
C a3 GND 10.8
R a3 5505
R adder_8_0/fulladder_5/a_85_7# 110
R adder_8_0/fulladder_5/a_77_7# 110
R adder_8_0/fulladder_5/a_45_7# 494
R adder_8_0/fulladder_5/a_29_7# 110
R adder_8_0/fulladder_5/a_n2_7# 504
R adder_8_0/fulladder_5/a_85_65# 281
R adder_8_0/fulladder_5/a_77_65# 281
R adder_8_0/fulladder_5/a_45_65# 838
R adder_8_0/fulladder_5/a_29_65# 281
R adder_8_0/fulladder_5/a_n2_65# 883
C adder_8_0/fulladder_5/a_69_7# GND 2.4
R adder_8_0/fulladder_5/a_69_7# 1250
C adder_8_0/fulladder_5/a_21_7# GND 5.8
R adder_8_0/fulladder_5/a_21_7# 2154
C adder_8_0/c_2_ GND 5.7
R adder_8_0/c_2_ 3139
C a2 GND 10.8
R a2 5505
R adder_8_0/fulladder_6/a_85_7# 110
R adder_8_0/fulladder_6/a_77_7# 110
R adder_8_0/fulladder_6/a_45_7# 494
R adder_8_0/fulladder_6/a_29_7# 110
R adder_8_0/fulladder_6/a_n2_7# 504
R adder_8_0/fulladder_6/a_85_65# 281
R adder_8_0/fulladder_6/a_77_65# 281
R adder_8_0/fulladder_6/a_45_65# 838
R adder_8_0/fulladder_6/a_29_65# 281
R adder_8_0/fulladder_6/a_n2_65# 883
C adder_8_0/fulladder_6/a_69_7# GND 2.4
R adder_8_0/fulladder_6/a_69_7# 1250
C adder_8_0/fulladder_6/a_21_7# GND 5.8
R adder_8_0/fulladder_6/a_21_7# 2154
C adder_8_0/c_1_ GND 5.7
R adder_8_0/c_1_ 3139
C a1 GND 10.9
R a1 5505
R adder_8_0/fulladder_7/a_85_7# 110
R adder_8_0/fulladder_7/a_77_7# 110
R adder_8_0/fulladder_7/a_45_7# 494
R adder_8_0/fulladder_7/a_29_7# 110
R adder_8_0/fulladder_7/a_n2_7# 504
R adder_8_0/fulladder_7/a_85_65# 281
R adder_8_0/fulladder_7/a_77_65# 281
R adder_8_0/fulladder_7/a_45_65# 838
R adder_8_0/fulladder_7/a_29_65# 281
R adder_8_0/fulladder_7/a_n2_65# 883
C adder_8_0/fulladder_7/a_69_7# GND 2.4
R adder_8_0/fulladder_7/a_69_7# 1250
C adder_8_0/fulladder_7/a_21_7# GND 5.8
R adder_8_0/fulladder_7/a_21_7# 2154
C a0 GND 11.5
R a0 5506
C mux3_1x_8_0/mux3_dp_1x_7/s0 GND 33.4
R mux3_1x_8_0/mux3_dp_1x_7/s0 9475
C mux3_1x_8_0/mux3_dp_1x_7/s0b GND 34.5
R mux3_1x_8_0/mux3_dp_1x_7/s0b 11370
C mux3_1x_8_0/mux3_dp_1x_7/s1 GND 39.0
R mux3_1x_8_0/mux3_dp_1x_7/s1 11502
C mux3_1x_8_0/mux3_dp_1x_7/s1b GND 35.3
R mux3_1x_8_0/mux3_dp_1x_7/s1b 11895
R mux3_1x_8_0/mux3_dp_1x_0/a_41_7# 164
R mux3_1x_8_0/mux3_dp_1x_0/a_20_7# 164
R mux3_1x_8_0/mux3_dp_1x_0/a_7_7# 164
R mux3_1x_8_0/mux3_dp_1x_0/a_0_7# 482
C result7 GND 8.4
R result7 1244
R mux3_1x_8_0/mux3_dp_1x_0/a_41_74# 316
C mux3_1x_8_0/mux3_dp_1x_0/a_33_7# GND 2.6
R mux3_1x_8_0/mux3_dp_1x_0/a_33_7# 1191
R mux3_1x_8_0/mux3_dp_1x_0/a_20_74# 316
R mux3_1x_8_0/mux3_dp_1x_0/a_7_74# 316
R mux3_1x_8_0/mux3_dp_1x_0/a_0_74# 668
C less GND 28.4
R less 9104
C adder_8_0/b_7_ GND 7.0
R adder_8_0/b_7_ 4907
C adder_8_0/s_7_ GND 3.1
R adder_8_0/s_7_ 1505
R mux3_1x_8_0/mux3_dp_1x_1/a_41_7# 164
R mux3_1x_8_0/mux3_dp_1x_1/a_20_7# 164
R mux3_1x_8_0/mux3_dp_1x_1/a_7_7# 164
R mux3_1x_8_0/mux3_dp_1x_1/a_0_7# 482
C result6 GND 9.2
R result6 1211
R mux3_1x_8_0/mux3_dp_1x_1/a_41_74# 316
C mux3_1x_8_0/mux3_dp_1x_1/a_33_7# GND 2.6
R mux3_1x_8_0/mux3_dp_1x_1/a_33_7# 1191
R mux3_1x_8_0/mux3_dp_1x_1/a_20_74# 316
R mux3_1x_8_0/mux3_dp_1x_1/a_7_74# 316
R mux3_1x_8_0/mux3_dp_1x_1/a_0_74# 668
C adder_8_0/b_6_ GND 7.5
R adder_8_0/b_6_ 4906
C adder_8_0/s_6_ GND 4.1
R adder_8_0/s_6_ 1506
R mux3_1x_8_0/mux3_dp_1x_2/a_41_7# 164
R mux3_1x_8_0/mux3_dp_1x_2/a_20_7# 164
R mux3_1x_8_0/mux3_dp_1x_2/a_7_7# 164
R mux3_1x_8_0/mux3_dp_1x_2/a_0_7# 482
C result5 GND 11.6
R result5 1246
R mux3_1x_8_0/mux3_dp_1x_2/a_41_74# 316
C mux3_1x_8_0/mux3_dp_1x_2/a_33_7# GND 2.6
R mux3_1x_8_0/mux3_dp_1x_2/a_33_7# 1191
R mux3_1x_8_0/mux3_dp_1x_2/a_20_74# 316
R mux3_1x_8_0/mux3_dp_1x_2/a_7_74# 316
R mux3_1x_8_0/mux3_dp_1x_2/a_0_74# 668
C adder_8_0/b_5_ GND 7.2
R adder_8_0/b_5_ 4906
C adder_8_0/s_5_ GND 4.1
R adder_8_0/s_5_ 1506
R mux3_1x_8_0/mux3_dp_1x_3/a_41_7# 164
R mux3_1x_8_0/mux3_dp_1x_3/a_20_7# 164
R mux3_1x_8_0/mux3_dp_1x_3/a_7_7# 164
R mux3_1x_8_0/mux3_dp_1x_3/a_0_7# 482
C result4 GND 9.2
R result4 1211
R mux3_1x_8_0/mux3_dp_1x_3/a_41_74# 316
C mux3_1x_8_0/mux3_dp_1x_3/a_33_7# GND 2.6
R mux3_1x_8_0/mux3_dp_1x_3/a_33_7# 1191
R mux3_1x_8_0/mux3_dp_1x_3/a_20_74# 316
R mux3_1x_8_0/mux3_dp_1x_3/a_7_74# 316
R mux3_1x_8_0/mux3_dp_1x_3/a_0_74# 668
C adder_8_0/b_4_ GND 7.0
R adder_8_0/b_4_ 4907
C adder_8_0/s_4_ GND 4.1
R adder_8_0/s_4_ 1506
R mux3_1x_8_0/mux3_dp_1x_4/a_41_7# 164
R mux3_1x_8_0/mux3_dp_1x_4/a_20_7# 164
R mux3_1x_8_0/mux3_dp_1x_4/a_7_7# 164
R mux3_1x_8_0/mux3_dp_1x_4/a_0_7# 482
C result3 GND 11.1
R result3 1245
R mux3_1x_8_0/mux3_dp_1x_4/a_41_74# 316
C mux3_1x_8_0/mux3_dp_1x_4/a_33_7# GND 2.6
R mux3_1x_8_0/mux3_dp_1x_4/a_33_7# 1191
R mux3_1x_8_0/mux3_dp_1x_4/a_20_74# 316
R mux3_1x_8_0/mux3_dp_1x_4/a_7_74# 316
R mux3_1x_8_0/mux3_dp_1x_4/a_0_74# 668
C adder_8_0/b_3_ GND 7.0
R adder_8_0/b_3_ 4907
C adder_8_0/s_3_ GND 4.1
R adder_8_0/s_3_ 1506
R mux3_1x_8_0/mux3_dp_1x_5/a_41_7# 164
R mux3_1x_8_0/mux3_dp_1x_5/a_20_7# 164
R mux3_1x_8_0/mux3_dp_1x_5/a_7_7# 164
R mux3_1x_8_0/mux3_dp_1x_5/a_0_7# 482
C result2 GND 9.1
R result2 1211
R mux3_1x_8_0/mux3_dp_1x_5/a_41_74# 316
C mux3_1x_8_0/mux3_dp_1x_5/a_33_7# GND 2.6
R mux3_1x_8_0/mux3_dp_1x_5/a_33_7# 1191
R mux3_1x_8_0/mux3_dp_1x_5/a_20_74# 316
R mux3_1x_8_0/mux3_dp_1x_5/a_7_74# 316
R mux3_1x_8_0/mux3_dp_1x_5/a_0_74# 668
C adder_8_0/b_2_ GND 7.0
R adder_8_0/b_2_ 4907
C adder_8_0/s_2_ GND 4.1
R adder_8_0/s_2_ 1506
R mux3_1x_8_0/mux3_dp_1x_6/a_41_7# 164
R mux3_1x_8_0/mux3_dp_1x_6/a_20_7# 164
R mux3_1x_8_0/mux3_dp_1x_6/a_7_7# 164
R mux3_1x_8_0/mux3_dp_1x_6/a_0_7# 482
C result1 GND 11.1
R result1 1245
R mux3_1x_8_0/mux3_dp_1x_6/a_41_74# 316
C mux3_1x_8_0/mux3_dp_1x_6/a_33_7# GND 2.6
R mux3_1x_8_0/mux3_dp_1x_6/a_33_7# 1191
R mux3_1x_8_0/mux3_dp_1x_6/a_20_74# 316
R mux3_1x_8_0/mux3_dp_1x_6/a_7_74# 316
R mux3_1x_8_0/mux3_dp_1x_6/a_0_74# 668
C adder_8_0/b_1_ GND 7.0
R adder_8_0/b_1_ 4907
C adder_8_0/s_1_ GND 4.1
R adder_8_0/s_1_ 1506
R mux3_1x_8_0/mux3_dp_1x_7/a_41_7# 164
R mux3_1x_8_0/mux3_dp_1x_7/a_20_7# 164
R mux3_1x_8_0/mux3_dp_1x_7/a_7_7# 164
R mux3_1x_8_0/mux3_dp_1x_7/a_0_7# 482
C result0 GND 9.9
R result0 1211
R mux3_1x_8_0/mux3_dp_1x_7/a_41_74# 316
C mux3_1x_8_0/mux3_dp_1x_7/a_33_7# GND 2.6
R mux3_1x_8_0/mux3_dp_1x_7/a_33_7# 1191
R mux3_1x_8_0/mux3_dp_1x_7/a_20_74# 316
R mux3_1x_8_0/mux3_dp_1x_7/a_7_74# 316
R mux3_1x_8_0/mux3_dp_1x_7/a_0_74# 668
C muxy7 GND 7.0
R muxy7 4907
C adder_8_0/s_0_ GND 4.1
R adder_8_0/s_0_ 1506
C Vdd! GND 1218.6
R Vdd! 268585
C op2 GND 23.4
R op2 4851
C funct_1 GND 41.9
R funct_1 6273
C alu_ctl_0/INVX2_0/Y GND 27.9
R alu_ctl_0/INVX2_0/Y 2229
C alu_ctl_0/OAI21X1_2/C GND 14.3
R alu_ctl_0/OAI21X1_2/C 3285
R alu_ctl_0/AOI21X1_0/a_12_6# 548
R alu_ctl_0/AOI21X1_0/a_2_54# 1765
C alu_op_0 GND 41.6
R alu_op_0 4314
C alu_ctl_0/INVX2_4/Y GND 7.6
R alu_ctl_0/INVX2_4/Y 2276
C op1 GND 18.7
R op1 3119
C alu_ctl_0/INVX2_1/A GND 23.0
R alu_ctl_0/INVX2_1/A 3628
R Gnd! 197884
C op0 GND 13.7
R op0 2007
R alu_ctl_0/OAI21X1_0/a_2_6# 800
R alu_ctl_0/OAI21X1_0/a_9_54# 1403
C alu_ctl_0/NAND3X1_2/Y GND 5.0
R alu_ctl_0/NAND3X1_2/Y 2556
C alu_op_1 GND 43.6
R alu_op_1 5441
R alu_ctl_0/OAI21X1_1/a_2_6# 800
R alu_ctl_0/OAI21X1_1/a_9_54# 1403
C alu_ctl_0/INVX2_2/Y GND 26.6
R alu_ctl_0/INVX2_2/Y 3327
C alu_ctl_0/INVX2_3/A GND 25.1
R alu_ctl_0/INVX2_3/A 3912
R alu_ctl_0/XOR2X1_0/a_35_6# 548
R alu_ctl_0/XOR2X1_0/a_18_6# 548
R alu_ctl_0/XOR2X1_0/a_35_54# 1403
C alu_ctl_0/XOR2X1_0/Y GND 7.5
R alu_ctl_0/XOR2X1_0/Y 1638
R alu_ctl_0/XOR2X1_0/a_18_54# 1403
C alu_ctl_0/XOR2X1_0/a_2_6# GND 3.5
R alu_ctl_0/XOR2X1_0/a_2_6# 2264
C alu_ctl_0/XOR2X1_0/a_13_43# GND 3.1
R alu_ctl_0/XOR2X1_0/a_13_43# 2220
C funct_2 GND 28.3
R funct_2 6535
C alu_ctl_0/INVX2_6/Y GND 6.5
R alu_ctl_0/INVX2_6/Y 2243
R alu_ctl_0/OAI21X1_2/a_2_6# 800
R alu_ctl_0/OAI21X1_2/a_9_54# 1403
C alu_ctl_0/OR2X1_0/Y GND 7.0
R alu_ctl_0/OR2X1_0/Y 1658
R alu_ctl_0/NAND2X1_0/a_9_6# 548
C alu_ctl_0/OAI21X1_2/B GND 6.0
R alu_ctl_0/OAI21X1_2/B 1730
C alu_ctl_0/INVX2_3/Y GND 9.6
R alu_ctl_0/INVX2_3/Y 3281
R alu_ctl_0/OAI21X1_3/a_2_6# 800
R alu_ctl_0/OAI21X1_3/a_9_54# 1403
R alu_ctl_0/OR2X1_0/a_9_54# 1403
C alu_ctl_0/OR2X1_0/a_2_54# GND 2.5
R alu_ctl_0/OR2X1_0/a_2_54# 2027
C funct_0 GND 42.3
R funct_0 6450
R alu_ctl_0/NAND2X1_1/a_9_6# 548
C alu_ctl_0/OAI21X1_7/B GND 10.9
R alu_ctl_0/OAI21X1_7/B 1731
R alu_ctl_0/AND2X2_0/a_9_6# 548
C alu_ctl_0/AND2X2_0/Y GND 13.1
R alu_ctl_0/AND2X2_0/Y 2260
C alu_ctl_0/AND2X2_0/a_2_6# GND 2.2
R alu_ctl_0/AND2X2_0/a_2_6# 1705
C funct_3 GND 20.9
R funct_3 2127
R alu_ctl_0/NAND3X1_0/a_14_6# 822
R alu_ctl_0/NAND3X1_0/a_9_6# 822
C alu_ctl_0/INVX2_5/Y GND 19.7
R alu_ctl_0/INVX2_5/Y 4431
R alu_ctl_0/OAI21X1_4/a_2_6# 800
C alu_ctl_0/NAND2X1_5/B GND 9.2
R alu_ctl_0/NAND2X1_5/B 2167
R alu_ctl_0/OAI21X1_4/a_9_54# 1403
C alu_ctl_0/NAND3X1_0/Y GND 9.6
R alu_ctl_0/NAND3X1_0/Y 3638
R alu_ctl_0/NAND2X1_2/a_9_6# 548
C alu_ctl_0/OAI21X1_7/A GND 9.2
R alu_ctl_0/OAI21X1_7/A 1754
R alu_ctl_0/NAND3X1_1/a_14_6# 822
R alu_ctl_0/NAND3X1_1/a_9_6# 822
C alu_ctl_0/NOR2X1_0/Y GND 4.6
R alu_ctl_0/NOR2X1_0/Y 1996
C funct_4 GND 13.7
R funct_4 1021
R alu_ctl_0/OAI21X1_5/a_2_6# 800
R alu_ctl_0/OAI21X1_5/a_9_54# 1403
C alu_ctl_0/INVX2_6/A GND 4.6
R alu_ctl_0/INVX2_6/A 2132
R alu_ctl_0/NAND2X1_3/a_9_6# 548
R alu_ctl_0/NAND3X1_2/a_14_6# 822
R alu_ctl_0/NAND3X1_2/a_9_6# 822
C alu_ctl_0/NOR2X1_0/A GND 13.9
R alu_ctl_0/NOR2X1_0/A 2761
R alu_ctl_0/NAND2X1_4/a_9_6# 548
R alu_ctl_0/OAI21X1_6/a_2_6# 800
R alu_ctl_0/OAI21X1_6/a_9_54# 1403
R alu_ctl_0/NAND2X1_5/a_9_6# 548
C alu_ctl_0/OAI21X1_6/C GND 3.9
R alu_ctl_0/OAI21X1_6/C 1717
C alu_ctl_0/NOR2X1_2/Y GND 13.6
R alu_ctl_0/NOR2X1_2/Y 4182
R alu_ctl_0/OAI21X1_7/a_2_6# 800
R alu_ctl_0/OAI21X1_7/a_9_54# 1403
R alu_ctl_0/NOR2X1_0/a_9_54# 1403
R alu_ctl_0/NOR2X1_1/a_9_54# 1403
R alu_ctl_0/NAND2X1_6/a_9_6# 548
C funct_5 GND 7.2
R funct_5 1050
C alu_ctl_0/NOR2X1_1/Y GND 4.8
R alu_ctl_0/NOR2X1_1/Y 1995
R alu_ctl_0/NOR2X1_2/a_9_54# 1403
C alu_ctl_0/NOR2X1_0/B GND 8.8
R alu_ctl_0/NOR2X1_0/B 2788
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        