magic
tech scmos
timestamp 1489863398
<< nwell >>
rect -6 40 50 96
<< ntransistor >>
rect 10 7 12 19
rect 15 7 17 19
rect 23 7 25 19
rect 28 7 30 19
rect 36 7 38 34
<< ptransistor >>
rect 10 65 12 83
rect 15 65 17 83
rect 23 65 25 83
rect 28 65 30 83
rect 36 46 38 83
<< ndiffusion >>
rect 31 32 36 34
rect 5 17 10 19
rect 9 8 10 17
rect 5 7 10 8
rect 12 7 15 19
rect 17 17 23 19
rect 17 8 18 17
rect 22 8 23 17
rect 17 7 23 8
rect 25 7 28 19
rect 30 8 31 19
rect 35 8 36 32
rect 30 7 36 8
rect 38 32 43 34
rect 38 8 39 32
rect 38 7 43 8
<< pdiffusion >>
rect 5 81 10 83
rect 9 67 10 81
rect 5 65 10 67
rect 12 65 15 83
rect 17 81 23 83
rect 17 67 18 81
rect 22 67 23 81
rect 17 65 23 67
rect 25 65 28 83
rect 30 81 36 83
rect 30 65 31 81
rect 35 52 36 81
rect 31 51 36 52
rect 33 46 36 51
rect 38 81 43 83
rect 38 47 39 81
rect 38 46 43 47
<< ndcontact >>
rect 5 8 9 17
rect 18 8 22 17
rect 31 8 35 32
rect 39 8 43 32
<< pdcontact >>
rect 5 67 9 81
rect 18 67 22 81
rect 31 52 35 81
rect 39 47 43 81
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
rect 40 -2 44 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
rect 32 88 36 92
rect 40 88 44 92
<< polysilicon >>
rect 10 83 12 85
rect 15 83 17 85
rect 23 83 25 85
rect 28 83 30 85
rect 36 83 38 85
rect 10 64 12 65
rect 2 62 12 64
rect 2 50 4 62
rect 15 59 17 65
rect 9 57 17 59
rect 9 50 11 57
rect 23 54 25 65
rect 18 53 25 54
rect 21 52 25 53
rect 2 6 4 46
rect 18 42 20 49
rect 28 48 30 65
rect 29 46 30 48
rect 10 40 20 42
rect 10 26 12 40
rect 27 33 29 44
rect 36 41 38 46
rect 37 37 38 41
rect 36 34 38 37
rect 27 31 30 33
rect 10 24 17 26
rect 10 19 12 21
rect 15 19 17 24
rect 20 22 22 30
rect 20 20 25 22
rect 23 19 25 20
rect 28 19 30 31
rect 10 6 12 7
rect 2 4 12 6
rect 15 5 17 7
rect 23 5 25 7
rect 28 5 30 7
rect 36 5 38 7
<< polycontact >>
rect 0 46 4 50
rect 8 46 12 50
rect 17 49 21 53
rect 25 44 29 48
rect 18 30 22 34
rect 33 37 37 41
<< metal1 >>
rect -2 92 46 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 32 92
rect 36 88 40 92
rect 44 88 46 92
rect -2 86 46 88
rect 5 81 9 86
rect 5 65 9 67
rect 18 81 22 83
rect 18 66 22 67
rect 20 62 22 66
rect 31 81 35 86
rect 18 55 24 59
rect 18 53 22 55
rect 31 51 35 52
rect 39 81 43 83
rect 8 34 12 46
rect 29 44 32 48
rect 43 47 44 50
rect 39 46 44 47
rect 40 42 44 46
rect 20 37 33 41
rect 40 34 44 38
rect 8 30 18 34
rect 31 32 35 34
rect 5 17 9 19
rect 20 17 22 19
rect 5 4 9 8
rect 18 7 22 8
rect 31 4 35 8
rect 39 32 44 34
rect 43 30 44 32
rect 39 7 43 8
rect -2 2 46 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 40 2
rect 44 -2 46 2
rect -2 -4 46 -2
<< m2contact >>
rect 16 62 20 66
rect 24 55 28 59
rect 0 46 4 50
rect 8 46 12 50
rect 32 44 36 48
rect 16 37 20 41
rect 40 38 44 42
rect 16 17 20 19
rect 16 15 18 17
rect 18 15 20 17
<< metal2 >>
rect 16 41 20 62
rect 16 19 20 37
<< labels >>
rlabel m2contact 2 48 2 48 1 d1
rlabel m2contact 10 48 10 48 1 sb
rlabel m2contact 26 57 26 57 1 s
rlabel m2contact 34 46 34 46 1 d0
rlabel m2contact 42 40 42 40 1 y
<< end >>
