magic
tech scmos
timestamp 1494266977
<< m2contact >>
rect -2 -2 2 2
<< end >>
