magic
tech scmos
timestamp 1484419411
<< nwell >>
rect -8 40 128 96
<< ntransistor >>
rect 3 7 5 15
rect 11 7 13 15
rect 19 7 21 15
rect 27 7 29 15
rect 35 7 37 15
rect 43 7 45 15
rect 51 7 53 15
rect 59 7 61 15
rect 67 7 69 15
rect 75 7 77 15
rect 83 7 85 15
rect 91 7 93 15
rect 99 7 101 15
rect 115 7 117 15
<< ptransistor >>
rect 3 65 5 81
rect 11 65 13 81
rect 19 65 21 81
rect 27 65 29 81
rect 35 65 37 81
rect 43 65 45 81
rect 51 65 53 81
rect 59 65 61 81
rect 67 65 69 81
rect 75 65 77 81
rect 83 65 85 81
rect 91 65 93 81
rect 99 65 101 81
rect 115 65 117 81
<< ndiffusion >>
rect 2 7 3 15
rect 5 7 6 15
rect 10 7 11 15
rect 13 7 14 15
rect 18 7 19 15
rect 21 7 22 15
rect 26 7 27 15
rect 29 7 35 15
rect 37 7 38 15
rect 42 7 43 15
rect 45 7 46 15
rect 50 7 51 15
rect 53 7 54 15
rect 58 7 59 15
rect 61 7 62 15
rect 66 7 67 15
rect 69 7 70 15
rect 74 7 75 15
rect 77 7 83 15
rect 85 7 91 15
rect 93 7 94 15
rect 98 7 99 15
rect 101 7 102 15
rect 114 7 115 15
rect 117 7 118 15
<< pdiffusion >>
rect -2 80 3 81
rect 2 66 3 80
rect -2 65 3 66
rect 5 72 6 81
rect 10 72 11 81
rect 5 65 11 72
rect 13 80 19 81
rect 13 66 14 80
rect 18 66 19 80
rect 13 65 19 66
rect 21 80 27 81
rect 21 67 22 80
rect 26 67 27 80
rect 21 65 27 67
rect 29 65 35 81
rect 37 80 43 81
rect 37 66 38 80
rect 42 66 43 80
rect 37 65 43 66
rect 45 80 51 81
rect 45 66 46 80
rect 50 66 51 80
rect 45 65 51 66
rect 53 72 54 81
rect 58 72 59 81
rect 53 65 59 72
rect 61 80 67 81
rect 61 66 62 80
rect 66 66 67 80
rect 61 65 67 66
rect 69 80 75 81
rect 69 67 70 80
rect 74 67 75 80
rect 69 65 75 67
rect 77 65 83 81
rect 85 65 91 81
rect 93 80 99 81
rect 93 66 94 80
rect 98 66 99 80
rect 93 65 99 66
rect 101 80 106 81
rect 101 67 102 80
rect 101 65 106 67
rect 110 80 115 81
rect 114 66 115 80
rect 110 65 115 66
rect 117 80 122 81
rect 117 66 118 80
rect 117 65 122 66
<< ndcontact >>
rect -2 7 2 15
rect 6 7 10 15
rect 14 7 18 15
rect 22 7 26 15
rect 38 7 42 15
rect 46 7 50 15
rect 54 7 58 15
rect 62 7 66 15
rect 70 7 74 15
rect 94 7 98 15
rect 102 7 106 15
rect 110 7 114 15
rect 118 7 122 15
<< pdcontact >>
rect -2 66 2 80
rect 6 72 10 81
rect 14 66 18 80
rect 22 67 26 80
rect 38 66 42 80
rect 46 66 50 80
rect 54 72 58 81
rect 62 66 66 80
rect 70 67 74 80
rect 94 66 98 80
rect 102 67 106 80
rect 110 66 114 80
rect 118 66 122 80
<< psubstratepcontact >>
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
<< nsubstratencontact >>
rect -2 88 2 92
rect 6 88 10 92
rect 14 88 18 92
rect 22 88 26 92
rect 30 88 34 92
rect 38 88 42 92
rect 46 88 50 92
rect 54 88 58 92
rect 62 88 66 92
rect 70 88 74 92
rect 78 88 82 92
rect 86 88 90 92
rect 94 88 98 92
rect 102 88 106 92
rect 110 88 114 92
rect 118 88 122 92
<< polysilicon >>
rect 3 81 5 83
rect 11 81 13 83
rect 19 81 21 83
rect 27 81 29 83
rect 35 81 37 83
rect 43 81 45 83
rect 51 81 53 83
rect 59 81 61 83
rect 67 81 69 83
rect 75 81 77 83
rect 83 81 85 83
rect 91 81 93 83
rect 99 81 101 83
rect 115 81 117 83
rect 3 36 5 65
rect 11 43 13 65
rect 19 51 21 65
rect 3 15 5 32
rect 11 15 13 39
rect 19 15 21 47
rect 27 43 29 65
rect 27 15 29 39
rect 35 36 37 65
rect 43 36 45 65
rect 51 43 53 65
rect 59 51 61 65
rect 35 15 37 32
rect 43 15 45 32
rect 51 15 53 39
rect 59 15 61 47
rect 67 29 69 65
rect 75 51 77 65
rect 67 15 69 25
rect 75 15 77 47
rect 83 43 85 65
rect 83 15 85 39
rect 91 36 93 65
rect 91 15 93 32
rect 99 22 101 65
rect 115 29 117 65
rect 99 15 101 18
rect 115 15 117 25
rect 3 5 5 7
rect 11 5 13 7
rect 19 5 21 7
rect 27 5 29 7
rect 35 5 37 7
rect 43 5 45 7
rect 51 5 53 7
rect 59 5 61 7
rect 67 5 69 7
rect 75 5 77 7
rect 83 5 85 7
rect 91 5 93 7
rect 99 5 101 7
rect 115 5 117 7
<< polycontact >>
rect 18 47 22 51
rect 10 39 14 43
rect 2 32 6 36
rect 26 39 30 43
rect 58 47 62 51
rect 50 39 54 43
rect 34 32 38 36
rect 42 32 46 36
rect 74 47 78 51
rect 66 25 70 29
rect 82 39 86 43
rect 90 32 94 36
rect 114 25 118 29
rect 98 18 102 22
<< metal1 >>
rect -4 92 124 94
rect -4 88 -2 92
rect 2 88 6 92
rect 10 88 14 92
rect 18 88 22 92
rect 26 88 30 92
rect 34 88 38 92
rect 42 88 46 92
rect 50 88 54 92
rect 58 88 62 92
rect 66 88 70 92
rect 74 88 78 92
rect 82 88 86 92
rect 90 88 94 92
rect 98 88 102 92
rect 106 88 110 92
rect 114 88 118 92
rect 122 88 124 92
rect -4 86 124 88
rect 6 81 10 86
rect -2 80 2 81
rect 14 80 18 81
rect 2 66 14 69
rect -2 65 18 66
rect 22 80 26 81
rect 38 80 42 86
rect 54 81 58 86
rect 38 65 42 66
rect 46 80 50 81
rect 62 80 66 81
rect 50 66 62 69
rect 46 65 66 66
rect 70 80 74 81
rect 94 80 98 86
rect 94 65 98 66
rect 102 80 106 81
rect 110 80 114 86
rect 110 65 114 66
rect 118 80 122 81
rect 118 59 122 66
rect 18 55 118 59
rect 22 47 58 51
rect 62 47 74 51
rect 14 39 26 43
rect 30 39 50 43
rect 54 39 82 43
rect 6 32 34 36
rect 38 32 42 36
rect 46 32 90 36
rect 26 25 66 29
rect 70 25 114 29
rect -2 18 18 22
rect -2 15 2 18
rect 14 15 18 18
rect 22 15 26 25
rect 46 18 66 22
rect 46 15 50 18
rect 62 15 66 18
rect 74 18 98 22
rect 70 15 74 18
rect 6 4 10 7
rect 38 4 42 7
rect 54 4 58 7
rect 94 4 98 7
rect 110 4 114 7
rect -4 2 124 4
rect -4 -2 -2 2
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 124 2
rect -4 -4 124 -2
<< m2contact >>
rect 22 67 26 69
rect 22 65 26 67
rect 70 67 74 69
rect 70 65 74 67
rect 102 67 106 69
rect 102 65 106 67
rect 14 55 18 59
rect 118 55 122 59
rect 14 47 18 51
rect 6 39 10 43
rect -2 32 2 36
rect 22 25 26 29
rect 70 18 74 22
rect 102 11 106 15
rect 118 11 122 15
<< metal2 >>
rect 22 29 26 65
rect 70 22 74 65
rect 102 15 106 65
rect 118 15 122 55
<< labels >>
rlabel m2contact 0 34 0 34 1 a
rlabel m2contact 8 41 8 41 1 b
rlabel m2contact 16 49 16 49 1 c
rlabel m2contact 16 57 16 57 1 cout
rlabel m2contact 104 13 104 13 1 s
rlabel metal1 4 89 4 89 1 Vdd!
rlabel metal1 4 -1 4 -1 1 Gnd!
<< end >>
