magic
tech scmos
timestamp 1484533619
<< ntransistor >>
rect 26 7 28 11
rect 56 7 58 11
<< ndiffusion >>
rect 25 7 26 11
rect 28 7 29 11
rect 55 7 56 11
rect 58 7 59 11
<< ndcontact >>
rect 21 7 25 11
rect 29 7 33 11
rect 51 7 55 11
rect 59 7 63 11
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
rect 40 -2 44 2
rect 48 -2 52 2
rect 56 -2 60 2
rect 64 -2 68 2
<< polysilicon >>
rect 24 14 26 18
rect 26 11 28 14
rect 56 11 58 14
rect 26 5 28 7
rect 56 5 58 7
<< polycontact >>
rect 26 14 30 18
rect 55 14 60 18
<< metal1 >>
rect 40 11 44 18
rect 33 7 44 11
rect 63 7 64 11
rect 21 4 25 7
rect 51 4 55 7
rect -2 2 70 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 40 2
rect 44 -2 48 2
rect 52 -2 56 2
rect 60 -2 64 2
rect 68 -2 70 2
rect -2 -4 70 -2
<< m2contact >>
rect 40 18 44 22
rect 24 14 26 18
rect 26 14 28 18
rect 56 14 60 18
rect 64 7 68 11
<< metal2 >>
rect 39 22 45 23
rect 39 18 40 22
rect 44 18 45 22
rect 39 17 45 18
rect 55 14 56 18
rect 63 12 69 13
rect 63 7 64 12
rect 68 7 69 12
<< m3contact >>
rect 40 18 44 22
rect 64 11 68 12
rect 64 8 68 11
<< metal3 >>
rect 39 22 45 23
rect 39 18 40 22
rect 44 18 45 22
rect 39 17 45 18
rect 63 12 69 13
rect 63 8 64 12
rect 68 8 69 12
rect 63 7 69 8
<< labels >>
rlabel m2contact 26 16 26 16 1 read1
rlabel m3contact 42 20 42 20 5 r1
rlabel m3contact 66 10 66 10 7 r2
rlabel m2contact 58 16 58 16 1 read2
<< end >>
