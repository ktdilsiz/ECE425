magic
tech scmos
timestamp 1488314249
<< error_s >>
rect 84 100 92 101
<< nwell >>
rect 80 97 84 101
<< metal1 >>
rect 22 860 30 868
rect 22 770 30 778
rect 22 750 30 758
rect 22 660 30 668
rect 22 640 30 648
rect 22 550 30 558
rect 22 530 30 538
rect 22 440 30 448
rect 22 420 30 428
rect 22 330 30 338
rect 22 310 30 318
rect 22 220 30 228
rect 22 200 30 208
rect 22 110 30 118
rect 22 90 30 98
rect 22 0 30 8
<< m2contact >>
rect 352 763 356 767
<< metal2 >>
rect 184 926 188 927
rect 48 837 52 838
rect 32 824 33 827
rect 32 812 36 824
rect 40 806 44 816
rect 48 812 52 833
rect 144 837 148 838
rect 144 830 148 833
rect 184 833 188 922
rect 273 876 277 926
rect 296 922 300 938
rect 328 922 332 929
rect 56 819 60 820
rect 56 815 57 819
rect 56 812 60 815
rect 0 670 4 711
rect 16 690 20 776
rect 48 727 52 728
rect 32 714 33 717
rect 32 702 36 714
rect 40 696 44 706
rect 48 702 52 723
rect 56 709 60 710
rect 56 705 57 709
rect 56 702 60 705
rect 48 617 52 618
rect 32 604 33 607
rect 32 592 36 604
rect 40 586 44 596
rect 48 592 52 613
rect 56 599 60 600
rect 56 595 57 599
rect 56 592 60 595
rect 0 450 4 491
rect 23 474 27 556
rect 48 507 52 508
rect 32 494 33 497
rect 32 482 36 494
rect 40 476 44 486
rect 48 482 52 503
rect 56 489 60 490
rect 56 485 57 489
rect 56 482 60 485
rect 48 397 52 398
rect 32 384 33 387
rect 32 372 36 384
rect 8 367 12 371
rect 40 366 44 376
rect 48 372 52 393
rect 56 379 60 380
rect 56 375 57 379
rect 56 372 60 375
rect 0 230 4 271
rect 16 250 20 336
rect 48 287 52 288
rect 32 274 33 277
rect 32 262 36 274
rect 40 256 44 266
rect 48 262 52 283
rect 56 269 60 270
rect 56 265 57 269
rect 56 262 60 265
rect 48 177 52 178
rect 32 168 36 169
rect 32 152 36 164
rect 40 146 44 156
rect 48 152 52 173
rect 56 159 60 160
rect 56 155 57 159
rect 56 152 60 155
rect 0 10 4 51
rect 16 30 20 116
rect 80 101 84 812
rect 48 67 52 68
rect 32 54 33 57
rect 32 42 36 54
rect 40 36 44 46
rect 48 42 52 63
rect 56 49 60 50
rect 56 45 57 49
rect 56 42 60 45
rect 80 38 84 97
rect 88 321 92 812
rect 112 806 116 812
rect 112 696 116 702
rect 112 586 116 592
rect 120 541 124 827
rect 160 811 164 813
rect 112 476 116 482
rect 112 366 116 372
rect 88 38 92 317
rect 112 256 116 262
rect 112 146 116 152
rect 96 53 100 54
rect 120 53 124 537
rect 136 761 140 811
rect 168 806 172 824
rect 312 817 316 826
rect 304 789 308 817
rect 112 36 116 42
rect 136 37 140 757
rect 144 727 148 728
rect 144 720 148 723
rect 160 701 164 703
rect 168 696 172 714
rect 312 707 316 716
rect 304 679 308 707
rect 144 617 148 618
rect 144 610 148 613
rect 160 591 164 593
rect 168 586 172 604
rect 312 597 316 606
rect 304 569 308 597
rect 144 507 148 508
rect 144 500 148 503
rect 160 481 164 483
rect 168 476 172 494
rect 312 487 316 496
rect 304 459 308 487
rect 144 397 148 398
rect 144 390 148 393
rect 160 371 164 373
rect 168 366 172 384
rect 312 377 316 386
rect 304 349 308 377
rect 144 287 148 288
rect 144 280 148 283
rect 160 261 164 263
rect 168 256 172 274
rect 312 267 316 276
rect 304 239 308 267
rect 144 177 148 178
rect 144 170 148 173
rect 160 151 164 153
rect 168 146 172 164
rect 312 157 316 166
rect 304 129 308 157
rect 144 67 148 68
rect 144 60 148 63
rect 279 58 283 106
rect 160 41 164 43
rect 168 36 172 54
rect 328 56 332 872
rect 352 767 356 826
rect 368 780 372 816
rect 352 104 356 763
rect 379 761 383 763
rect 368 670 372 706
rect 379 702 383 757
rect 368 560 372 596
rect 379 492 383 537
rect 368 450 372 486
rect 368 340 372 376
rect 379 272 383 317
rect 368 230 372 266
rect 368 120 372 156
rect 389 110 393 917
rect 379 62 383 97
rect 184 51 188 52
rect 312 47 316 56
rect 304 19 308 47
rect 368 10 372 46
<< m3contact >>
rect 296 938 300 942
rect 691 938 695 942
rect 184 922 188 926
rect 265 922 269 926
rect 48 833 52 837
rect 33 824 37 828
rect 144 833 148 837
rect 328 929 332 933
rect 395 929 399 933
rect 389 917 393 921
rect 273 872 277 876
rect 328 872 332 876
rect 184 829 188 833
rect 95 824 100 828
rect 57 815 61 819
rect 64 815 68 819
rect 40 802 44 806
rect 16 776 20 780
rect 48 723 52 727
rect 33 714 37 718
rect 57 705 61 709
rect 64 705 68 709
rect 40 692 44 696
rect 0 666 4 670
rect 48 613 52 617
rect 33 604 37 608
rect 57 595 61 599
rect 64 595 68 599
rect 40 582 44 586
rect 23 556 27 560
rect 48 503 52 507
rect 33 494 37 498
rect 16 470 20 474
rect 23 470 27 474
rect 57 485 61 489
rect 64 485 68 489
rect 40 472 44 476
rect 0 446 4 450
rect 48 393 52 397
rect 33 384 37 388
rect 57 375 61 379
rect 64 375 68 379
rect 40 362 44 366
rect 16 336 20 340
rect 48 283 52 287
rect 33 274 37 278
rect 57 265 61 269
rect 64 265 68 269
rect 40 252 44 256
rect 0 226 4 230
rect 48 173 52 177
rect 32 164 36 168
rect 57 155 61 159
rect 64 155 68 159
rect 40 142 44 146
rect 16 116 20 120
rect 80 97 84 101
rect 48 63 52 67
rect 33 54 37 58
rect 57 45 61 49
rect 64 45 68 49
rect 112 802 116 806
rect 95 714 100 718
rect 112 692 116 696
rect 95 604 100 608
rect 112 582 116 586
rect 168 824 172 828
rect 160 813 164 817
rect 120 537 124 541
rect 95 494 100 498
rect 112 472 116 476
rect 95 384 100 388
rect 112 362 116 366
rect 88 317 92 321
rect 95 274 100 278
rect 112 252 116 256
rect 95 164 100 168
rect 112 142 116 146
rect 95 54 100 58
rect 176 813 180 817
rect 312 813 316 817
rect 272 785 276 789
rect 304 785 308 789
rect 136 757 140 761
rect 40 32 44 36
rect 144 723 148 727
rect 168 714 172 718
rect 160 703 164 707
rect 176 703 180 707
rect 312 703 316 707
rect 272 675 276 679
rect 304 675 308 679
rect 144 613 148 617
rect 168 604 172 608
rect 160 593 164 597
rect 176 593 180 597
rect 312 593 316 597
rect 272 565 276 569
rect 304 565 308 569
rect 144 503 148 507
rect 168 494 172 498
rect 160 483 164 487
rect 176 483 180 487
rect 312 483 316 487
rect 272 455 276 459
rect 304 455 308 459
rect 144 393 148 397
rect 168 384 172 388
rect 160 373 164 377
rect 176 373 180 377
rect 312 373 316 377
rect 272 345 276 349
rect 304 345 308 349
rect 144 283 148 287
rect 168 274 172 278
rect 160 263 164 267
rect 176 263 180 267
rect 312 263 316 267
rect 272 235 276 239
rect 304 235 308 239
rect 144 173 148 177
rect 168 164 172 168
rect 160 153 164 157
rect 176 153 180 157
rect 312 153 316 157
rect 272 125 276 129
rect 304 125 308 129
rect 279 106 283 110
rect 144 63 148 67
rect 168 54 172 58
rect 160 43 164 47
rect 184 52 188 56
rect 279 54 283 58
rect 368 776 372 780
rect 379 757 383 761
rect 379 698 383 702
rect 368 666 372 670
rect 368 556 372 560
rect 379 537 383 541
rect 379 488 383 492
rect 368 446 372 450
rect 368 336 372 340
rect 379 317 383 321
rect 379 268 383 272
rect 368 226 372 230
rect 368 116 372 120
rect 389 106 393 110
rect 379 97 383 101
rect 379 58 383 62
rect 328 52 332 56
rect 352 52 356 56
rect 176 43 180 47
rect 112 32 116 36
rect 312 43 316 47
rect 272 15 276 19
rect 304 15 308 19
rect 0 6 4 10
rect 368 6 372 10
<< metal3 >>
rect 295 942 697 943
rect 295 938 296 942
rect 300 938 691 942
rect 695 938 697 942
rect 295 937 697 938
rect 327 933 400 934
rect 327 929 328 933
rect 332 929 395 933
rect 399 929 400 933
rect 327 928 400 929
rect 183 926 270 927
rect 183 922 184 926
rect 188 922 265 926
rect 269 922 270 926
rect 183 921 270 922
rect 388 921 394 922
rect 388 917 389 921
rect 393 917 394 921
rect 388 916 394 917
rect 272 876 333 877
rect 272 872 273 876
rect 277 872 328 876
rect 332 872 333 876
rect 272 871 333 872
rect 47 837 149 838
rect 47 833 48 837
rect 52 833 144 837
rect 148 833 149 837
rect 47 832 149 833
rect 183 833 189 834
rect 183 829 184 833
rect 188 829 189 833
rect 32 828 173 829
rect 183 828 189 829
rect 32 824 33 828
rect 37 824 95 828
rect 100 824 168 828
rect 172 824 173 828
rect 32 823 173 824
rect 56 819 69 820
rect 56 815 57 819
rect 61 815 64 819
rect 68 815 69 819
rect 56 814 69 815
rect 159 817 317 818
rect 159 813 160 817
rect 164 813 176 817
rect 180 813 312 817
rect 316 813 317 817
rect 159 812 317 813
rect 39 806 117 807
rect 39 802 40 806
rect 44 802 112 806
rect 116 802 117 806
rect 39 801 117 802
rect 271 789 309 790
rect 271 785 272 789
rect 276 785 304 789
rect 308 785 309 789
rect 271 784 309 785
rect -2 780 373 781
rect -2 776 16 780
rect 20 776 368 780
rect 372 776 373 780
rect -2 775 373 776
rect 135 761 384 762
rect 135 757 136 761
rect 140 757 379 761
rect 383 757 384 761
rect 135 756 384 757
rect 47 727 149 728
rect 47 723 48 727
rect 52 723 144 727
rect 148 723 149 727
rect 47 722 149 723
rect 32 718 173 719
rect 32 714 33 718
rect 37 714 95 718
rect 100 714 168 718
rect 172 714 173 718
rect 32 713 173 714
rect 56 709 69 710
rect 56 705 57 709
rect 61 705 64 709
rect 68 705 69 709
rect 56 704 69 705
rect 159 707 317 708
rect 159 703 160 707
rect 164 703 176 707
rect 180 703 312 707
rect 316 703 317 707
rect 159 702 317 703
rect 378 702 384 703
rect 378 698 379 702
rect 383 698 384 702
rect 378 697 384 698
rect 39 696 117 697
rect 39 692 40 696
rect 44 692 112 696
rect 116 692 117 696
rect 39 691 117 692
rect 271 679 309 680
rect 271 675 272 679
rect 276 675 304 679
rect 308 675 309 679
rect 271 674 309 675
rect -2 670 373 671
rect -2 666 0 670
rect 4 666 368 670
rect 372 666 373 670
rect -2 665 373 666
rect 47 617 149 618
rect 47 613 48 617
rect 52 613 144 617
rect 148 613 149 617
rect 47 612 149 613
rect 32 608 173 609
rect 32 604 33 608
rect 37 604 95 608
rect 100 604 168 608
rect 172 604 173 608
rect 32 603 173 604
rect 56 599 69 600
rect 56 595 57 599
rect 61 595 64 599
rect 68 595 69 599
rect 56 594 69 595
rect 159 597 317 598
rect 159 593 160 597
rect 164 593 176 597
rect 180 593 312 597
rect 316 593 317 597
rect 159 592 317 593
rect 39 586 117 587
rect 39 582 40 586
rect 44 582 112 586
rect 116 582 117 586
rect 39 581 117 582
rect 271 569 309 570
rect 271 565 272 569
rect 276 565 304 569
rect 308 565 309 569
rect 271 564 309 565
rect -2 560 373 561
rect -2 556 23 560
rect 27 556 368 560
rect 372 556 373 560
rect -2 555 373 556
rect 119 541 384 542
rect 119 537 120 541
rect 124 537 379 541
rect 383 537 384 541
rect 119 536 384 537
rect 47 507 149 508
rect 47 503 48 507
rect 52 503 144 507
rect 148 503 149 507
rect 47 502 149 503
rect 32 498 173 499
rect 32 494 33 498
rect 37 494 95 498
rect 100 494 168 498
rect 172 494 173 498
rect 32 493 173 494
rect 378 492 384 493
rect 56 489 69 490
rect 56 485 57 489
rect 61 485 64 489
rect 68 485 69 489
rect 378 488 379 492
rect 383 488 384 492
rect 56 484 69 485
rect 159 487 317 488
rect 378 487 384 488
rect 159 483 160 487
rect 164 483 176 487
rect 180 483 312 487
rect 316 483 317 487
rect 159 482 317 483
rect 39 476 117 477
rect 15 474 28 475
rect 15 470 16 474
rect 20 470 23 474
rect 27 470 28 474
rect 39 472 40 476
rect 44 472 112 476
rect 116 472 117 476
rect 39 471 117 472
rect 15 469 28 470
rect 271 459 309 460
rect 271 455 272 459
rect 276 455 304 459
rect 308 455 309 459
rect 271 454 309 455
rect -2 450 373 451
rect -2 446 0 450
rect 4 446 368 450
rect 372 446 373 450
rect -2 445 373 446
rect 47 397 149 398
rect 47 393 48 397
rect 52 393 144 397
rect 148 393 149 397
rect 47 392 149 393
rect 32 388 173 389
rect 32 384 33 388
rect 37 384 95 388
rect 100 384 168 388
rect 172 384 173 388
rect 32 383 173 384
rect 56 379 69 380
rect 56 375 57 379
rect 61 375 64 379
rect 68 375 69 379
rect 56 374 69 375
rect 159 377 317 378
rect 159 373 160 377
rect 164 373 176 377
rect 180 373 312 377
rect 316 373 317 377
rect 159 372 317 373
rect 39 366 117 367
rect 39 362 40 366
rect 44 362 112 366
rect 116 362 117 366
rect 39 361 117 362
rect 271 349 309 350
rect 271 345 272 349
rect 276 345 304 349
rect 308 345 309 349
rect 271 344 309 345
rect -2 340 373 341
rect -2 336 16 340
rect 20 336 368 340
rect 372 336 373 340
rect -2 335 373 336
rect 87 321 384 322
rect 87 317 88 321
rect 92 317 379 321
rect 383 317 384 321
rect 87 316 384 317
rect 47 287 149 288
rect 47 283 48 287
rect 52 283 144 287
rect 148 283 149 287
rect 47 282 149 283
rect 32 278 173 279
rect 32 274 33 278
rect 37 274 95 278
rect 100 274 168 278
rect 172 274 173 278
rect 32 273 173 274
rect 378 272 384 273
rect 56 269 69 270
rect 56 265 57 269
rect 61 265 64 269
rect 68 265 69 269
rect 378 268 379 272
rect 383 268 384 272
rect 56 264 69 265
rect 159 267 317 268
rect 378 267 384 268
rect 159 263 160 267
rect 164 263 176 267
rect 180 263 312 267
rect 316 263 317 267
rect 159 262 317 263
rect 39 256 117 257
rect 39 252 40 256
rect 44 252 112 256
rect 116 252 117 256
rect 39 251 117 252
rect 271 239 309 240
rect 271 235 272 239
rect 276 235 304 239
rect 308 235 309 239
rect 271 234 309 235
rect -2 230 373 231
rect -2 226 0 230
rect 4 226 368 230
rect 372 226 373 230
rect -2 225 373 226
rect 47 177 149 178
rect 47 173 48 177
rect 52 173 144 177
rect 148 173 149 177
rect 47 172 149 173
rect 31 168 173 169
rect 31 164 32 168
rect 36 164 95 168
rect 100 164 168 168
rect 172 164 173 168
rect 31 163 173 164
rect 56 159 69 160
rect 56 155 57 159
rect 61 155 64 159
rect 68 155 69 159
rect 56 154 69 155
rect 159 157 317 158
rect 159 153 160 157
rect 164 153 176 157
rect 180 153 312 157
rect 316 153 317 157
rect 159 152 317 153
rect 39 146 117 147
rect 39 142 40 146
rect 44 142 112 146
rect 116 142 117 146
rect 39 141 117 142
rect 271 129 309 130
rect 271 125 272 129
rect 276 125 304 129
rect 308 125 309 129
rect 271 124 309 125
rect -2 120 373 121
rect -2 116 16 120
rect 20 116 368 120
rect 372 116 373 120
rect -2 115 373 116
rect 278 110 395 111
rect 278 106 279 110
rect 283 106 389 110
rect 393 106 395 110
rect 278 105 395 106
rect 79 101 384 102
rect 79 97 80 101
rect 84 97 379 101
rect 383 97 384 101
rect 79 96 384 97
rect 47 67 149 68
rect 47 63 48 67
rect 52 63 144 67
rect 148 63 149 67
rect 47 62 149 63
rect 378 62 384 63
rect 32 58 173 59
rect 32 54 33 58
rect 37 54 95 58
rect 100 54 168 58
rect 172 54 173 58
rect 32 53 173 54
rect 183 58 284 59
rect 183 56 279 58
rect 183 52 184 56
rect 188 54 279 56
rect 283 54 284 58
rect 378 58 379 62
rect 383 58 384 62
rect 378 57 384 58
rect 188 53 284 54
rect 327 56 357 57
rect 188 52 189 53
rect 183 51 189 52
rect 327 52 328 56
rect 332 52 352 56
rect 356 52 357 56
rect 327 51 357 52
rect 56 49 69 50
rect 56 45 57 49
rect 61 45 64 49
rect 68 45 69 49
rect 56 44 69 45
rect 159 47 317 48
rect 159 43 160 47
rect 164 43 176 47
rect 180 43 312 47
rect 316 43 317 47
rect 159 42 317 43
rect 39 36 117 37
rect 39 32 40 36
rect 44 32 112 36
rect 116 32 117 36
rect 39 31 117 32
rect 271 19 309 20
rect 271 15 272 19
rect 276 15 304 19
rect 308 15 309 19
rect 271 14 309 15
rect -2 10 373 11
rect -2 6 0 10
rect 4 6 368 10
rect 372 6 373 10
rect -2 5 373 6
use inv_1x  inv_1x_0
timestamp 1484418501
transform 1 0 265 0 1 884
box -6 -4 18 96
use yzdetect_8  yzdetect_8_0
timestamp 1484534894
transform 1 0 0 0 1 4
box -8 -4 28 756
use inv_1x_8  inv_1x_8_0
timestamp 1484534894
transform 1 0 32 0 1 4
box -6 -4 18 866
use inv_1x_8  inv_1x_8_1
timestamp 1484534894
transform 1 0 48 0 1 4
box -6 -4 18 866
use mux4_8_10space  mux4_8_10space_0
timestamp 1487099744
transform 1 0 58 0 1 0
box 0 0 112 870
use adder_8  adder_8_0
timestamp 1484427118
transform 1 0 168 0 1 4
box -6 -4 130 866
use mux3_1x_8  mux3_1x_8_0
timestamp 1484532969
transform 1 0 296 0 1 4
box -6 -4 82 976
use alu_ctl  alu_ctl_0
timestamp 1488311641
transform 1 0 378 0 1 0
box 0 0 400 980
<< labels >>
rlabel metal2 33 46 33 46 1 a0
rlabel metal2 49 46 49 46 1 b0
rlabel metal2 33 156 33 156 1 a1
rlabel metal2 49 156 49 156 1 b1
rlabel metal2 33 266 33 266 1 a2
rlabel metal2 49 266 49 266 1 b2
rlabel metal2 33 376 33 376 1 a3
rlabel metal2 49 376 49 376 1 b3
rlabel metal2 33 486 33 486 1 a4
rlabel metal2 49 486 49 486 1 b4
rlabel metal2 33 596 33 596 1 a5
rlabel metal3 -1 9 -1 9 1 result0
rlabel metal3 -1 119 -1 119 1 result1
rlabel metal3 -1 230 -1 230 1 result2
rlabel metal3 -1 340 -1 340 1 result3
rlabel metal3 -1 450 -1 450 1 result4
rlabel metal3 -1 560 -1 560 1 result5
rlabel metal3 -1 670 -1 670 1 result6
rlabel metal3 1 778 1 778 1 result7
rlabel m2contact 352 763 356 767 1 less
rlabel metal2 296 922 300 926 1 op0
rlabel metal2 328 922 332 926 1 op1
rlabel metal2 49 596 49 596 1 b5
rlabel metal2 33 706 33 706 1 a6
rlabel metal2 49 706 49 706 1 b6
rlabel metal2 33 816 33 816 1 a7
rlabel metal2 49 816 49 816 1 b7
rlabel metal2 9 370 9 370 1 zero
rlabel m3contact 161 44 161 44 1 muxy7
rlabel metal2 81 767 81 767 1 op6
rlabel metal2 89 767 89 767 1 op5
rlabel metal2 120 763 124 767 1 op4
rlabel metal2 136 763 140 767 1 op3
rlabel m3contact 98 56 98 56 1 mux4s1_0
rlabel metal2 146 61 146 61 1 mux4s0_0
rlabel m3contact 186 830 186 830 1 cout_adder_7
rlabel metal2 122 544 122 544 1 op4
rlabel metal2 90 325 90 325 1 op5
rlabel metal2 82 104 82 104 1 op6
rlabel metal2 186 52 186 52 1 op2
rlabel metal2 281 106 281 106 1 op2
<< end >>
