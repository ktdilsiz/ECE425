magic
tech scmos
timestamp 1484532969
<< metal1 >>
rect -2 966 38 974
rect -2 876 38 884
rect 12 868 24 872
rect 44 868 56 872
<< m2contact >>
rect 8 868 12 872
rect 24 868 28 872
rect 40 868 44 872
rect 56 868 60 872
<< metal2 >>
rect -1 902 5 903
rect -1 898 0 902
rect 4 898 5 902
rect -1 897 5 898
rect 0 49 4 897
rect 8 872 12 923
rect 24 903 28 921
rect 40 903 44 921
rect 23 902 29 903
rect 23 898 24 902
rect 28 898 29 902
rect 23 897 29 898
rect 38 902 44 903
rect 38 898 39 902
rect 43 898 44 902
rect 38 897 44 898
rect 47 902 53 903
rect 47 898 48 902
rect 52 898 53 902
rect 47 897 53 898
rect 24 49 28 868
rect 40 40 44 868
rect 48 49 52 897
rect 56 872 60 922
<< m3contact >>
rect 0 898 4 902
rect 24 898 28 902
rect 39 898 43 902
rect 48 898 52 902
<< metal3 >>
rect -1 902 29 903
rect -1 898 0 902
rect 4 898 24 902
rect 28 898 29 902
rect -1 897 29 898
rect 38 902 53 903
rect 38 898 39 902
rect 43 898 48 902
rect 52 898 53 902
rect 38 897 53 898
use invbuf_4x  invbuf_4x_0
timestamp 1484532969
transform 1 0 0 0 1 880
box -6 -4 34 96
use invbuf_4x  invbuf_4x_1
timestamp 1484532969
transform 1 0 32 0 1 880
box -6 -4 34 96
use mux3_dp_1x  mux3_dp_1x_0
timestamp 1484514831
transform 1 0 0 0 1 770
box -6 -4 82 96
use mux3_dp_1x  mux3_dp_1x_1
timestamp 1484514831
transform 1 0 0 0 1 660
box -6 -4 82 96
use mux3_dp_1x  mux3_dp_1x_2
timestamp 1484514831
transform 1 0 0 0 1 550
box -6 -4 82 96
use mux3_dp_1x  mux3_dp_1x_3
timestamp 1484514831
transform 1 0 0 0 1 440
box -6 -4 82 96
use mux3_dp_1x  mux3_dp_1x_4
timestamp 1484514831
transform 1 0 0 0 1 330
box -6 -4 82 96
use mux3_dp_1x  mux3_dp_1x_5
timestamp 1484514831
transform 1 0 0 0 1 220
box -6 -4 82 96
use mux3_dp_1x  mux3_dp_1x_6
timestamp 1484514831
transform 1 0 0 0 1 110
box -6 -4 82 96
use mux3_dp_1x  mux3_dp_1x_7
timestamp 1484514831
transform 1 0 0 0 1 0
box -6 -4 82 96
<< end >>
