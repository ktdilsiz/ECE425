magic
tech scmos
timestamp 1493662838
<< nwell >>
rect -6 40 147 96
<< ntransistor >>
rect 13 8 15 32
rect 21 14 23 32
rect 27 15 29 21
rect 35 15 37 21
rect 40 15 42 21
rect 61 8 63 14
rect 69 8 71 12
rect 76 8 78 12
rect 85 8 87 14
rect 93 8 95 14
rect 101 8 103 12
rect 108 8 110 12
rect 117 8 119 14
rect 133 8 135 15
<< ptransistor >>
rect 13 71 15 83
rect 18 71 20 83
rect 26 77 28 83
rect 31 77 33 83
rect 39 77 41 83
rect 61 77 63 83
rect 69 79 71 83
rect 76 79 78 83
rect 85 74 87 83
rect 93 77 95 83
rect 101 79 103 83
rect 108 79 110 83
rect 117 74 119 83
rect 133 73 135 83
<< ndiffusion >>
rect 12 8 13 32
rect 15 8 16 32
rect 20 14 21 32
rect 23 21 26 32
rect 23 15 27 21
rect 29 20 35 21
rect 29 16 30 20
rect 34 16 35 20
rect 29 15 35 16
rect 37 15 40 21
rect 42 20 47 21
rect 42 16 43 20
rect 42 15 47 16
rect 23 14 26 15
rect 60 8 61 14
rect 63 8 64 14
rect 80 13 85 14
rect 68 8 69 12
rect 71 8 76 12
rect 78 9 80 12
rect 84 9 85 13
rect 78 8 85 9
rect 87 8 88 14
rect 92 8 93 14
rect 95 8 96 14
rect 100 8 101 12
rect 103 8 108 12
rect 110 8 112 12
rect 116 8 117 14
rect 119 8 120 14
rect 132 8 133 15
rect 135 8 136 15
<< pdiffusion >>
rect 8 81 13 83
rect 12 72 13 81
rect 8 71 13 72
rect 15 71 18 83
rect 20 81 26 83
rect 20 72 21 81
rect 25 77 26 81
rect 28 77 31 83
rect 33 82 39 83
rect 33 78 34 82
rect 38 78 39 82
rect 33 77 39 78
rect 41 82 46 83
rect 41 78 42 82
rect 41 77 46 78
rect 56 82 61 83
rect 60 78 61 82
rect 56 77 61 78
rect 63 77 64 83
rect 68 79 69 83
rect 71 79 76 83
rect 78 79 80 83
rect 20 71 25 72
rect 84 74 85 83
rect 87 74 88 83
rect 92 77 93 83
rect 95 77 96 83
rect 100 79 101 83
rect 103 79 108 83
rect 110 79 112 83
rect 116 74 117 83
rect 119 74 120 83
rect 128 82 133 83
rect 132 73 133 82
rect 135 82 140 83
rect 135 73 136 82
<< ndcontact >>
rect 8 8 12 32
rect 16 8 20 32
rect 30 16 34 20
rect 43 16 47 20
rect 56 8 60 14
rect 64 8 68 14
rect 80 9 84 13
rect 88 8 92 14
rect 96 8 100 14
rect 112 8 116 14
rect 120 8 124 14
rect 128 8 132 15
rect 136 8 140 15
<< pdcontact >>
rect 8 72 12 81
rect 21 72 25 81
rect 34 78 38 82
rect 42 78 46 82
rect 56 78 60 82
rect 64 77 68 83
rect 80 74 84 83
rect 88 74 92 83
rect 96 77 100 83
rect 112 74 116 83
rect 120 74 124 83
rect 128 73 132 82
rect 136 73 140 82
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
rect 40 -2 44 2
rect 48 -2 52 2
rect 56 -2 60 2
rect 64 -2 68 2
rect 72 -2 76 2
rect 80 -2 84 2
rect 88 -2 92 2
rect 96 -2 100 2
rect 104 -2 108 2
rect 112 -2 116 2
rect 120 -2 124 2
rect 128 -2 132 2
rect 136 -2 140 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
rect 32 88 36 92
rect 40 88 44 92
rect 48 88 52 92
rect 56 88 60 92
rect 64 88 68 92
rect 72 88 76 92
rect 80 88 84 92
rect 88 88 92 92
rect 96 88 100 92
rect 104 88 108 92
rect 112 88 116 92
rect 120 88 124 92
rect 128 88 132 92
rect 136 88 140 92
<< polysilicon >>
rect 13 83 15 85
rect 18 83 20 85
rect 26 83 28 85
rect 31 83 33 85
rect 39 83 41 85
rect 61 83 63 85
rect 69 83 71 85
rect 76 83 78 85
rect 85 83 87 85
rect 93 83 95 85
rect 101 83 103 85
rect 108 83 110 85
rect 117 83 119 85
rect 133 83 135 85
rect 13 66 15 71
rect 14 63 15 66
rect 18 66 20 71
rect 18 64 23 66
rect 13 32 15 53
rect 21 47 23 64
rect 26 55 28 77
rect 31 61 33 77
rect 39 69 41 77
rect 39 67 46 69
rect 31 59 39 61
rect 26 53 34 55
rect 24 43 29 46
rect 21 32 23 35
rect 27 21 29 43
rect 32 36 34 53
rect 37 49 39 59
rect 44 57 46 67
rect 61 57 63 77
rect 69 74 71 79
rect 76 67 78 79
rect 76 63 77 67
rect 37 47 40 49
rect 61 45 63 53
rect 61 43 71 45
rect 32 34 49 36
rect 35 21 37 34
rect 40 26 41 30
rect 40 21 42 26
rect 21 12 23 14
rect 27 13 29 15
rect 35 13 37 15
rect 40 13 42 15
rect 61 14 63 17
rect 69 12 71 43
rect 76 12 78 63
rect 85 28 87 74
rect 93 57 95 77
rect 101 74 103 79
rect 108 67 110 79
rect 108 63 109 67
rect 96 53 103 55
rect 86 24 87 28
rect 85 14 87 24
rect 93 14 95 17
rect 101 12 103 53
rect 108 12 110 63
rect 117 37 119 74
rect 118 33 119 37
rect 117 14 119 33
rect 133 15 135 73
rect 13 6 15 8
rect 61 6 63 8
rect 69 6 71 8
rect 76 6 78 8
rect 85 6 87 8
rect 93 6 95 8
rect 101 6 103 8
rect 108 6 110 8
rect 117 6 119 8
rect 133 6 135 8
<< polycontact >>
rect 10 62 14 66
rect 12 53 16 57
rect 20 43 24 47
rect 19 35 23 39
rect 68 70 72 74
rect 77 63 81 67
rect 43 53 47 57
rect 60 53 64 57
rect 40 45 44 49
rect 49 33 53 37
rect 41 26 45 30
rect 60 17 64 21
rect 100 70 104 74
rect 109 63 113 67
rect 92 53 96 57
rect 82 24 86 28
rect 92 17 96 21
rect 129 41 133 45
rect 114 33 118 37
<< metal1 >>
rect -2 92 142 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 32 92
rect 36 88 40 92
rect 44 88 48 92
rect 52 88 56 92
rect 60 88 64 92
rect 68 88 72 92
rect 76 88 80 92
rect 84 88 88 92
rect 92 88 96 92
rect 100 88 104 92
rect 108 88 112 92
rect 116 88 120 92
rect 124 88 128 92
rect 132 88 136 92
rect 140 88 142 92
rect -2 86 142 88
rect 8 81 12 86
rect 8 71 12 72
rect 21 81 25 83
rect 34 82 38 86
rect 80 83 84 86
rect 112 83 116 86
rect 34 77 38 78
rect 42 82 46 83
rect 42 74 46 78
rect 25 72 32 74
rect 21 70 32 72
rect 36 71 46 74
rect 56 82 60 83
rect 56 71 60 78
rect 36 70 56 71
rect 42 67 56 70
rect 88 67 92 74
rect 120 67 124 74
rect 128 82 132 86
rect 136 82 140 83
rect 4 62 10 66
rect 14 62 40 64
rect 10 60 40 62
rect 81 63 88 67
rect 113 63 124 67
rect 20 53 43 57
rect 64 53 80 57
rect 96 53 112 57
rect 40 39 44 45
rect 52 43 72 47
rect 120 45 124 63
rect 124 41 129 45
rect 136 42 140 73
rect 12 35 19 39
rect 23 35 44 39
rect 53 33 96 37
rect 100 33 114 37
rect 30 22 32 26
rect 68 24 82 28
rect 30 20 34 22
rect 104 21 108 25
rect 30 15 34 16
rect 43 20 47 21
rect 64 17 72 21
rect 96 17 108 21
rect 43 12 47 16
rect 136 15 140 38
rect 20 8 47 12
rect 80 13 84 14
rect 8 4 12 8
rect 80 4 84 9
rect 112 4 116 8
rect 128 4 132 8
rect -2 2 142 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 40 2
rect 44 -2 48 2
rect 52 -2 56 2
rect 60 -2 64 2
rect 68 -2 72 2
rect 76 -2 80 2
rect 84 -2 88 2
rect 92 -2 96 2
rect 100 -2 104 2
rect 108 -2 112 2
rect 116 -2 120 2
rect 124 -2 128 2
rect 132 -2 136 2
rect 140 -2 142 2
rect -2 -4 142 -2
<< m2contact >>
rect 32 70 36 74
rect 64 77 68 81
rect 96 77 100 81
rect 56 67 60 71
rect 72 70 76 74
rect 104 70 108 74
rect 0 62 4 66
rect 40 60 44 64
rect 88 63 92 67
rect 16 53 20 57
rect 80 53 84 57
rect 112 53 116 57
rect 24 43 28 47
rect 48 43 52 47
rect 72 43 76 47
rect 120 41 124 45
rect 8 35 12 39
rect 136 38 140 42
rect 96 33 100 37
rect 40 26 41 30
rect 41 26 44 30
rect 32 22 36 26
rect 64 24 68 28
rect 104 25 108 29
rect 72 17 76 21
rect 56 10 60 14
rect 64 10 68 14
rect 88 10 92 14
rect 96 10 100 14
rect 120 10 124 14
<< metal2 >>
rect 32 26 36 70
rect 40 30 44 60
rect 56 14 60 67
rect 64 28 68 77
rect 64 14 68 24
rect 72 47 76 70
rect 72 21 76 43
rect 88 14 92 63
rect 96 37 100 77
rect 96 14 100 33
rect 104 29 108 70
rect 120 14 124 41
<< labels >>
rlabel m2contact 2 64 2 64 1 enb
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel m2contact 10 37 10 37 1 en
rlabel m2contact 26 45 26 45 1 d
rlabel m2contact 50 45 50 45 1 ph2
rlabel m2contact 106 27 106 27 1 ph1
rlabel m2contact 138 40 138 40 1 q
rlabel m2contact 114 55 114 55 1 phi1b
rlabel m2contact 82 55 82 55 1 phi2b
rlabel metal1 6 0 6 0 1 Gnd!
rlabel m2contact 18 55 18 55 1 resetb
rlabel metal2 90 39 90 39 1 master
rlabel metal2 98 39 98 39 1 slave
<< end >>
