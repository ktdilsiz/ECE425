magic
tech scmos
timestamp 1490727624
<< m2contact >>
rect -7 -7 7 7
<< end >>
