magic
tech scmos
timestamp 1485570478
<< nwell >>
rect 26 40 146 96
<< ntransistor >>
rect 37 8 39 32
rect 45 8 47 14
rect 61 8 63 14
rect 69 8 71 12
rect 76 8 78 12
rect 85 8 87 14
rect 93 8 95 14
rect 101 8 103 12
rect 108 8 110 12
rect 117 8 119 14
rect 133 7 135 34
<< ptransistor >>
rect 37 71 39 83
rect 45 77 47 83
rect 61 77 63 83
rect 69 79 71 83
rect 76 79 78 83
rect 85 74 87 83
rect 93 77 95 83
rect 101 79 103 83
rect 108 79 110 83
rect 117 74 119 83
rect 133 46 135 83
<< ndiffusion >>
rect 36 8 37 32
rect 39 8 40 32
rect 44 8 45 14
rect 47 8 48 14
rect 60 8 61 14
rect 63 8 64 14
rect 80 13 85 14
rect 68 8 69 12
rect 71 8 76 12
rect 78 9 80 12
rect 84 9 85 13
rect 78 8 85 9
rect 87 8 88 14
rect 92 8 93 14
rect 95 8 96 14
rect 128 32 133 34
rect 112 13 117 14
rect 100 8 101 12
rect 103 8 108 12
rect 110 9 112 12
rect 116 9 117 13
rect 110 8 117 9
rect 119 8 120 14
rect 132 8 133 32
rect 128 7 133 8
rect 135 32 140 34
rect 135 8 136 32
rect 135 7 140 8
<< pdiffusion >>
rect 32 81 37 83
rect 36 72 37 81
rect 32 71 37 72
rect 39 81 45 83
rect 39 72 40 81
rect 44 77 45 81
rect 47 82 52 83
rect 47 78 48 82
rect 47 77 52 78
rect 56 82 61 83
rect 60 78 61 82
rect 56 77 61 78
rect 63 77 64 83
rect 68 79 69 83
rect 71 79 76 83
rect 78 79 80 83
rect 39 71 44 72
rect 84 74 85 83
rect 87 74 88 83
rect 92 77 93 83
rect 95 77 96 83
rect 100 79 101 83
rect 103 79 108 83
rect 110 79 112 83
rect 116 74 117 83
rect 119 74 120 83
rect 128 81 133 83
rect 132 47 133 81
rect 128 46 133 47
rect 135 81 140 83
rect 135 47 136 81
rect 135 46 140 47
<< ndcontact >>
rect 32 8 36 32
rect 40 8 44 32
rect 48 8 52 14
rect 56 8 60 14
rect 64 8 68 14
rect 80 9 84 13
rect 88 8 92 14
rect 96 8 100 14
rect 112 9 116 13
rect 120 8 124 14
rect 128 8 132 32
rect 136 8 140 32
<< pdcontact >>
rect 32 72 36 81
rect 40 72 44 81
rect 48 78 52 82
rect 56 78 60 82
rect 64 77 68 83
rect 80 74 84 83
rect 88 74 92 83
rect 96 77 100 83
rect 112 74 116 83
rect 120 74 124 83
rect 128 47 132 81
rect 136 47 140 81
<< psubstratepcontact >>
rect 32 -2 36 2
rect 40 -2 44 2
rect 48 -2 52 2
rect 56 -2 60 2
rect 64 -2 68 2
rect 72 -2 76 2
rect 80 -2 84 2
rect 88 -2 92 2
rect 96 -2 100 2
rect 104 -2 108 2
rect 112 -2 116 2
rect 120 -2 124 2
rect 128 -2 132 2
rect 136 -2 140 2
<< nsubstratencontact >>
rect 32 88 36 92
rect 40 88 44 92
rect 48 88 52 92
rect 56 88 60 92
rect 64 88 68 92
rect 72 88 76 92
rect 80 88 84 92
rect 88 88 92 92
rect 96 88 100 92
rect 104 88 108 92
rect 112 88 116 92
rect 120 88 124 92
rect 128 88 132 92
rect 136 88 140 92
<< polysilicon >>
rect 37 83 39 85
rect 45 83 47 85
rect 61 83 63 85
rect 69 83 71 85
rect 76 83 78 85
rect 85 83 87 85
rect 93 83 95 85
rect 101 83 103 85
rect 108 83 110 85
rect 117 83 119 85
rect 133 83 135 85
rect 37 63 39 71
rect 45 69 47 77
rect 45 67 54 69
rect 37 61 47 63
rect 37 32 39 53
rect 45 47 47 61
rect 52 57 54 67
rect 61 57 63 77
rect 69 74 71 79
rect 76 67 78 79
rect 76 63 77 67
rect 61 45 63 53
rect 61 43 71 45
rect 45 14 47 43
rect 61 14 63 17
rect 69 12 71 43
rect 76 12 78 63
rect 85 28 87 74
rect 93 57 95 77
rect 101 74 103 79
rect 108 67 110 79
rect 108 63 109 67
rect 96 53 103 55
rect 86 24 87 28
rect 85 14 87 24
rect 93 14 95 17
rect 101 12 103 53
rect 108 12 110 63
rect 117 36 119 74
rect 118 32 119 36
rect 133 34 135 46
rect 117 14 119 32
rect 37 6 39 8
rect 45 6 47 8
rect 61 6 63 8
rect 69 6 71 8
rect 76 6 78 8
rect 85 6 87 8
rect 93 6 95 8
rect 101 6 103 8
rect 108 6 110 8
rect 117 6 119 8
rect 133 5 135 7
<< polycontact >>
rect 36 53 40 57
rect 68 70 72 74
rect 77 63 81 67
rect 52 53 56 57
rect 60 53 64 57
rect 44 43 48 47
rect 60 17 64 21
rect 100 70 104 74
rect 109 63 113 67
rect 92 53 96 57
rect 82 24 86 28
rect 92 17 96 21
rect 129 39 133 43
rect 114 32 118 36
<< metal1 >>
rect 30 92 142 94
rect 30 88 32 92
rect 36 88 40 92
rect 44 88 48 92
rect 52 88 56 92
rect 60 88 64 92
rect 68 88 72 92
rect 76 88 80 92
rect 84 88 88 92
rect 92 88 96 92
rect 100 88 104 92
rect 108 88 112 92
rect 116 88 120 92
rect 124 88 128 92
rect 132 88 136 92
rect 140 88 142 92
rect 30 86 142 88
rect 32 81 36 86
rect 40 81 44 83
rect 32 71 36 72
rect 39 72 40 75
rect 48 82 52 86
rect 80 83 84 86
rect 112 83 116 86
rect 48 77 52 78
rect 56 82 60 83
rect 56 74 60 78
rect 44 72 56 74
rect 39 70 56 72
rect 88 67 92 74
rect 120 67 124 74
rect 81 63 88 67
rect 113 63 124 67
rect 44 53 52 57
rect 64 53 80 57
rect 96 53 112 57
rect 120 43 124 63
rect 128 81 132 86
rect 128 46 132 47
rect 136 81 140 83
rect 136 43 140 47
rect 124 39 129 43
rect 48 30 56 34
rect 100 33 114 36
rect 96 32 114 33
rect 128 32 132 34
rect 48 14 52 30
rect 68 24 82 28
rect 104 21 108 25
rect 64 17 72 21
rect 96 17 108 21
rect 80 13 84 14
rect 32 4 36 8
rect 80 4 84 9
rect 112 13 116 14
rect 112 4 116 9
rect 128 4 132 8
rect 136 32 140 39
rect 136 7 140 8
rect 30 2 142 4
rect 30 -2 32 2
rect 36 -2 40 2
rect 44 -2 48 2
rect 52 -2 56 2
rect 60 -2 64 2
rect 68 -2 72 2
rect 76 -2 80 2
rect 84 -2 88 2
rect 92 -2 96 2
rect 100 -2 104 2
rect 108 -2 112 2
rect 116 -2 120 2
rect 124 -2 128 2
rect 132 -2 136 2
rect 140 -2 142 2
rect 30 -4 142 -2
<< m2contact >>
rect 64 77 68 81
rect 96 77 100 81
rect 56 70 60 74
rect 72 70 76 74
rect 104 70 108 74
rect 88 63 92 67
rect 40 53 44 57
rect 80 53 84 57
rect 112 53 116 57
rect 48 43 52 47
rect 72 43 76 47
rect 120 39 124 43
rect 136 39 140 43
rect 56 30 60 34
rect 96 33 100 37
rect 64 24 68 28
rect 104 25 108 29
rect 72 17 76 21
rect 56 10 60 14
rect 64 10 68 14
rect 88 10 92 14
rect 96 10 100 14
rect 120 10 124 14
<< metal2 >>
rect 56 34 60 70
rect 56 14 60 30
rect 64 28 68 77
rect 64 14 68 24
rect 72 47 76 70
rect 72 21 76 43
rect 88 14 92 63
rect 96 37 100 77
rect 96 14 100 33
rect 104 29 108 70
rect 120 14 124 39
<< labels >>
rlabel metal1 31 -1 31 -1 2 Gnd!
rlabel metal1 31 90 31 90 3 Vdd!
rlabel m2contact 50 45 50 45 1 d
rlabel m2contact 42 55 42 55 1 resetb
rlabel m2contact 74 45 74 45 1 ph2
rlabel m2contact 82 55 82 55 1 ph2b
rlabel m2contact 114 55 114 55 1 ph1b
rlabel m2contact 98 35 98 35 1 ph1
rlabel m2contact 138 41 138 41 1 q
<< end >>
