magic
tech scmos
timestamp 1484411102
<< nwell >>
rect -6 40 26 96
<< ntransistor >>
rect 5 7 7 15
rect 13 7 15 15
<< ptransistor >>
rect 5 67 7 83
rect 10 67 12 83
<< ndiffusion >>
rect 0 13 5 15
rect 4 9 5 13
rect 0 7 5 9
rect 7 13 13 15
rect 7 9 8 13
rect 12 9 13 13
rect 7 7 13 9
rect 15 13 20 15
rect 15 9 16 13
rect 15 7 20 9
<< pdiffusion >>
rect 0 82 5 83
rect 4 68 5 82
rect 0 67 5 68
rect 7 67 10 83
rect 12 82 17 83
rect 12 68 13 82
rect 12 67 17 68
<< ndcontact >>
rect 0 9 4 13
rect 8 9 12 13
rect 16 9 20 13
<< pdcontact >>
rect 0 68 4 82
rect 13 68 17 82
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
<< polysilicon >>
rect 5 83 7 85
rect 10 83 12 85
rect 5 47 7 67
rect 1 43 2 47
rect 6 43 7 47
rect 5 15 7 43
rect 10 44 12 67
rect 10 42 15 44
rect 13 15 15 42
rect 5 5 7 7
rect 13 5 15 7
<< polycontact >>
rect 2 43 6 47
rect 15 26 19 30
<< metal1 >>
rect -2 92 22 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 22 92
rect -2 86 22 88
rect 0 82 4 86
rect 0 67 4 68
rect 13 82 17 83
rect 13 37 17 68
rect 12 33 17 37
rect 0 13 4 15
rect 0 4 4 9
rect 8 13 12 33
rect 8 7 12 9
rect 16 13 20 15
rect 16 4 20 9
rect -2 2 22 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 22 2
rect -2 -4 22 -2
<< m2contact >>
rect 0 43 2 47
rect 2 43 4 47
rect 8 33 12 37
rect 16 26 19 30
rect 19 26 20 30
<< labels >>
rlabel m2contact 2 45 2 45 1 a
rlabel m2contact 10 35 10 35 1 y
rlabel m2contact 18 28 18 28 1 b
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel metal1 -1 0 -1 0 3 Gnd!
<< end >>
