magic
tech scmos
timestamp 1490643393
<< nwell >>
rect -48 16 14 76
<< ntransistor >>
rect -37 -9 -35 6
rect -29 -9 -27 6
rect -13 -9 -11 6
rect -5 -9 -3 6
<< ptransistor >>
rect -37 27 -35 57
rect -29 27 -27 57
rect -13 27 -11 57
rect -5 27 -3 57
<< ndiffusion >>
rect -42 -3 -37 6
rect -38 -7 -37 -3
rect -42 -9 -37 -7
rect -35 -3 -29 6
rect -35 -7 -34 -3
rect -30 -7 -29 -3
rect -35 -9 -29 -7
rect -27 -3 -22 6
rect -27 -7 -26 -3
rect -27 -9 -22 -7
rect -18 -3 -13 6
rect -14 -7 -13 -3
rect -18 -9 -13 -7
rect -11 -3 -5 6
rect -11 -7 -10 -3
rect -6 -7 -5 -3
rect -11 -9 -5 -7
rect -3 -3 2 6
rect -3 -7 -2 -3
rect -3 -9 2 -7
<< pdiffusion >>
rect -38 27 -37 57
rect -35 27 -34 57
rect -30 27 -29 57
rect -27 27 -26 57
rect -14 27 -13 57
rect -11 27 -10 57
rect -6 27 -5 57
rect -3 27 -2 57
<< ndcontact >>
rect -42 -7 -38 -3
rect -34 -7 -30 -3
rect -26 -7 -22 -3
rect -18 -7 -14 -3
rect -10 -7 -6 -3
rect -2 -7 2 -3
<< pdcontact >>
rect -42 27 -38 57
rect -34 27 -30 57
rect -26 27 -22 57
rect -18 27 -14 57
rect -10 27 -6 57
rect -2 27 2 57
<< psubstratepcontact >>
rect -42 -18 -38 -14
rect -34 -18 -30 -14
rect -26 -18 -22 -14
rect -18 -18 -14 -14
rect -10 -18 -6 -14
rect -2 -18 2 -14
rect 6 -18 10 -14
<< nsubstratencontact >>
rect -42 69 -38 73
rect -34 69 -30 73
rect -26 69 -22 73
rect -18 69 -14 73
rect -10 69 -6 73
rect -2 69 2 73
rect 6 69 10 73
<< polysilicon >>
rect -37 57 -35 59
rect -29 57 -27 59
rect -13 57 -11 59
rect -5 57 -3 59
rect -37 23 -35 27
rect -43 19 -42 23
rect -38 19 -35 23
rect -37 16 -35 19
rect -29 16 -27 27
rect -37 14 -27 16
rect -37 6 -35 14
rect -29 6 -27 14
rect -13 13 -11 27
rect -5 13 -3 27
rect -13 11 7 13
rect -13 6 -11 11
rect -5 6 -3 11
rect 5 6 7 11
rect -37 -11 -35 -9
rect -29 -11 -27 -9
rect -13 -11 -11 -9
rect -5 -11 -3 -9
<< polycontact >>
rect -42 19 -38 23
rect 5 2 9 6
<< metal1 >>
rect -46 73 12 75
rect -46 69 -42 73
rect -38 69 -34 73
rect -30 69 -26 73
rect -22 69 -18 73
rect -14 69 -10 73
rect -6 69 -2 73
rect 2 69 6 73
rect 10 69 12 73
rect -46 67 12 69
rect -42 57 -38 67
rect -26 57 -22 67
rect -10 60 9 64
rect -10 57 -6 60
rect -34 23 -30 27
rect -18 23 -14 27
rect -2 23 2 27
rect -34 19 2 23
rect 5 37 9 60
rect 5 13 9 33
rect -34 9 9 13
rect -42 -3 -38 6
rect -42 -12 -38 -7
rect -34 -3 -30 9
rect -34 -9 -30 -7
rect -26 -3 -22 6
rect -26 -12 -22 -7
rect -18 -3 -14 6
rect -18 -12 -14 -7
rect -10 -3 -6 9
rect -10 -9 -6 -7
rect -2 -3 2 6
rect -2 -12 2 -7
rect -46 -14 12 -12
rect -46 -18 -42 -14
rect -38 -18 -34 -14
rect -30 -18 -26 -14
rect -22 -18 -18 -14
rect -14 -18 -10 -14
rect -6 -18 -2 -14
rect 2 -18 6 -14
rect 10 -18 12 -14
rect -46 -20 12 -18
<< m2contact >>
rect -44 19 -42 23
rect -42 19 -40 23
rect 5 33 9 37
rect 6 2 9 6
rect 9 2 10 6
<< labels >>
rlabel metal1 -43 -16 -43 -16 3 Gnd!
rlabel m2contact 7 35 7 35 1 y
rlabel metal1 -43 71 -43 71 3 Vdd!
rlabel m2contact 8 4 8 4 1 b
rlabel m2contact -42 21 -42 21 1 a
<< end >>
