magic
tech scmos
timestamp 1484418501
<< nwell >>
rect -6 40 18 96
<< ntransistor >>
rect 5 7 7 14
<< ptransistor >>
rect 5 73 7 83
<< ndiffusion >>
rect 0 12 5 14
rect 4 8 5 12
rect 0 7 5 8
rect 7 12 12 14
rect 7 8 8 12
rect 7 7 12 8
<< pdiffusion >>
rect 0 82 5 83
rect 4 73 5 82
rect 7 82 12 83
rect 7 73 8 82
<< ndcontact >>
rect 0 8 4 12
rect 8 8 12 12
<< pdcontact >>
rect 0 73 4 82
rect 8 73 12 82
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
<< polysilicon >>
rect 5 83 7 85
rect 5 14 7 73
rect 5 5 7 7
<< polycontact >>
rect 1 38 5 42
<< metal1 >>
rect -2 92 14 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 14 92
rect -2 86 14 88
rect 0 82 4 86
rect 8 82 12 83
rect 8 42 12 73
rect 0 12 4 14
rect 0 4 4 8
rect 8 12 12 38
rect 8 7 12 8
rect -2 2 14 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 14 2
rect -2 -4 14 -2
<< m2contact >>
rect 0 38 1 42
rect 1 38 4 42
rect 8 38 12 42
<< labels >>
rlabel m2contact 1 40 1 40 1 a
rlabel m2contact 10 40 10 40 1 y
rlabel metal1 -1 0 -1 0 3 Gnd!
rlabel metal1 -1 90 -1 90 3 Vdd!
<< end >>
