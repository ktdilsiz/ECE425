magic
tech scmos
timestamp 1487689792
<< nwell >>
rect -6 40 34 96
<< ntransistor >>
rect 5 7 7 31
rect 10 7 12 31
rect 15 7 17 31
<< ptransistor >>
rect 5 63 7 83
rect 13 63 15 83
rect 21 63 23 83
<< ndiffusion >>
rect 4 7 5 31
rect 7 7 10 31
rect 12 7 15 31
rect 17 7 18 31
<< pdiffusion >>
rect 0 82 5 83
rect 4 63 5 82
rect 7 82 13 83
rect 7 63 8 82
rect 12 63 13 82
rect 15 82 21 83
rect 15 63 16 82
rect 20 63 21 82
rect 23 82 28 83
rect 23 63 24 82
<< ndcontact >>
rect 0 7 4 31
rect 18 7 22 31
<< pdcontact >>
rect 0 63 4 82
rect 8 63 12 82
rect 16 63 20 82
rect 24 63 28 82
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
<< polysilicon >>
rect 5 83 7 85
rect 13 83 15 85
rect 21 83 23 85
rect 5 62 7 63
rect 13 62 15 63
rect 1 60 7 62
rect 10 60 15 62
rect 1 47 3 60
rect 10 47 12 60
rect 21 58 23 63
rect 18 56 23 58
rect 18 47 20 56
rect 1 34 3 43
rect 1 32 7 34
rect 5 31 7 32
rect 10 31 12 43
rect 18 34 20 43
rect 15 32 20 34
rect 15 31 17 32
rect 5 5 7 7
rect 10 5 12 7
rect 15 5 17 7
<< polycontact >>
rect 0 43 4 47
rect 8 43 12 47
rect 16 43 20 47
<< metal1 >>
rect -2 92 30 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 30 92
rect -2 86 30 88
rect 0 82 4 86
rect 8 82 12 83
rect 16 82 20 86
rect 24 82 28 83
rect 8 60 12 63
rect 24 60 28 63
rect 8 56 28 60
rect 24 47 28 56
rect 24 31 28 43
rect 22 27 28 31
rect 0 4 4 7
rect -2 2 30 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 30 2
rect -2 -4 30 -2
<< m2contact >>
rect 0 43 4 47
rect 8 43 12 47
rect 16 43 20 47
rect 24 43 28 47
<< labels >>
rlabel m2contact 2 45 2 45 1 a
rlabel m2contact 10 45 10 45 1 b
rlabel m2contact 18 45 18 45 1 c
rlabel m2contact 26 45 26 45 1 y
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel metal1 -1 0 -1 0 3 Gnd!
<< end >>
