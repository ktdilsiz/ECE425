magic
tech scmos
timestamp 1487714794
<< nwell >>
rect -6 40 42 96
<< ntransistor >>
rect 5 28 7 32
rect 10 28 12 32
rect 18 28 20 32
rect 21 17 25 19
<< ptransistor >>
rect 24 75 28 77
rect 5 59 7 63
rect 13 59 15 63
rect 21 59 23 63
<< ndiffusion >>
rect 4 28 5 32
rect 7 28 10 32
rect 12 28 13 32
rect 17 28 18 32
rect 20 28 21 32
rect 21 19 25 20
rect 21 16 25 17
<< pdiffusion >>
rect 24 77 28 78
rect 24 74 28 75
rect 4 59 5 63
rect 7 59 8 63
rect 12 59 13 63
rect 15 59 16 63
rect 20 59 21 63
rect 23 59 24 63
<< ndcontact >>
rect 0 28 4 32
rect 13 28 17 32
rect 21 28 25 32
rect 21 20 25 24
rect 21 12 25 16
<< pdcontact >>
rect 24 78 28 82
rect 24 70 28 74
rect 0 59 4 63
rect 8 59 12 63
rect 16 59 20 63
rect 24 59 28 63
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
rect 32 88 36 92
<< polysilicon >>
rect 22 75 24 77
rect 28 75 31 77
rect 5 63 7 65
rect 13 63 15 65
rect 21 63 23 65
rect 5 55 7 59
rect 13 55 15 59
rect 21 55 23 59
rect 0 53 7 55
rect 10 53 15 55
rect 18 53 23 55
rect 0 47 2 53
rect 10 47 12 53
rect 18 47 20 53
rect 0 37 2 43
rect 0 35 7 37
rect 5 32 7 35
rect 10 32 12 43
rect 18 32 20 43
rect 29 37 31 75
rect 5 26 7 28
rect 10 26 12 28
rect 18 26 20 28
rect 26 19 28 36
rect 19 17 21 19
rect 25 17 28 19
<< polycontact >>
rect 0 43 4 47
rect 8 43 12 47
rect 16 43 20 47
rect 25 36 29 40
<< metal1 >>
rect -2 92 38 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 32 92
rect 36 88 38 92
rect -2 86 38 88
rect 13 74 17 86
rect 28 78 32 82
rect 8 70 24 74
rect 8 63 12 70
rect 0 55 4 59
rect 16 55 20 59
rect 0 51 20 55
rect 24 40 28 59
rect 13 36 25 40
rect 13 32 17 36
rect 0 24 4 28
rect 21 24 25 28
rect 0 20 21 24
rect 7 4 11 20
rect 25 12 32 16
rect -2 2 38 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 38 2
rect -2 -4 38 -2
<< m2contact >>
rect 32 78 36 82
rect 0 43 4 47
rect 8 43 12 47
rect 16 43 20 47
rect 32 12 36 16
<< metal2 >>
rect 32 16 36 78
<< labels >>
rlabel m2contact 2 45 2 45 1 a
rlabel m2contact 10 45 10 45 1 b
rlabel m2contact 18 45 18 45 1 c
rlabel metal2 34 45 34 45 1 y
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel metal1 -1 0 -1 0 3 Gnd!
<< end >>
