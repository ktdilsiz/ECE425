magic
tech scmos
timestamp 1489946810
<< nwell >>
rect -6 40 42 96
<< ntransistor >>
rect 5 7 7 27
rect 10 7 12 27
rect 15 7 17 27
rect 20 7 22 27
<< ptransistor >>
rect 5 69 7 83
rect 13 69 15 83
rect 21 69 23 83
rect 29 69 31 83
<< ndiffusion >>
rect 0 26 5 27
rect 4 7 5 26
rect 7 7 10 27
rect 12 7 15 27
rect 17 7 20 27
rect 22 26 27 27
rect 22 7 23 26
<< pdiffusion >>
rect 4 69 5 83
rect 7 69 8 83
rect 12 69 13 83
rect 15 69 16 83
rect 20 69 21 83
rect 23 69 24 83
rect 28 69 29 83
rect 31 69 32 83
<< ndcontact >>
rect 0 7 4 26
rect 23 7 27 26
<< pdcontact >>
rect 0 69 4 83
rect 8 69 12 83
rect 16 69 20 83
rect 24 69 28 83
rect 32 69 36 83
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
rect 32 88 36 92
<< polysilicon >>
rect 5 83 7 85
rect 13 83 15 85
rect 21 83 23 85
rect 29 83 31 85
rect 5 60 7 69
rect 13 68 15 69
rect 0 58 7 60
rect 10 66 15 68
rect 0 55 4 58
rect 0 39 2 51
rect 0 37 7 39
rect 5 27 7 37
rect 10 27 12 66
rect 21 47 23 69
rect 15 43 16 47
rect 20 45 23 47
rect 15 27 17 43
rect 29 39 31 69
rect 20 37 31 39
rect 20 27 22 37
rect 5 5 7 7
rect 10 5 12 7
rect 15 5 17 7
rect 20 5 22 7
<< polycontact >>
rect 0 51 4 55
rect 6 43 10 47
rect 16 43 20 47
rect 31 43 35 47
<< metal1 >>
rect -2 92 38 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 32 92
rect 36 88 38 92
rect -2 86 38 88
rect 0 83 4 86
rect 16 83 20 86
rect 32 83 36 86
rect 8 58 12 69
rect 24 58 28 69
rect 8 57 28 58
rect 8 54 24 57
rect 23 53 24 54
rect 0 26 4 27
rect 23 26 27 53
rect 0 4 4 7
rect -2 2 38 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 38 2
rect -2 -4 38 -2
<< m2contact >>
rect 0 55 4 57
rect 0 53 4 55
rect 24 53 28 57
rect 8 43 10 47
rect 10 43 12 47
rect 16 43 20 47
rect 33 43 35 47
rect 35 43 37 47
<< metal2 >>
rect 31 43 33 47
<< labels >>
rlabel m2contact 35 45 35 45 1 d
rlabel m2contact 26 55 26 55 1 y
rlabel m2contact 18 45 18 45 1 c
rlabel m2contact 10 45 10 45 1 b
rlabel m2contact 2 55 2 55 1 a
<< end >>
