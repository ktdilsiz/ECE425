magic
tech scmos
timestamp 1484419186
<< nwell >>
rect -6 40 106 96
<< ntransistor >>
rect 11 7 13 13
rect 16 7 18 13
rect 24 7 26 13
rect 29 7 31 13
rect 37 7 39 13
rect 45 7 47 13
rect 53 7 55 13
rect 58 7 60 13
rect 66 7 68 13
rect 71 7 73 13
rect 93 7 95 14
<< ptransistor >>
rect 11 74 13 83
rect 16 74 18 83
rect 24 74 26 83
rect 29 74 31 83
rect 37 74 39 83
rect 45 74 47 83
rect 53 74 55 83
rect 58 74 60 83
rect 66 74 68 83
rect 71 74 73 83
rect 93 73 95 83
<< ndiffusion >>
rect 6 12 11 13
rect 10 8 11 12
rect 6 7 11 8
rect 13 7 16 13
rect 18 12 24 13
rect 18 8 19 12
rect 23 8 24 12
rect 18 7 24 8
rect 26 7 29 13
rect 31 12 37 13
rect 31 8 32 12
rect 36 8 37 12
rect 31 7 37 8
rect 39 12 45 13
rect 39 8 40 12
rect 44 8 45 12
rect 39 7 45 8
rect 47 12 53 13
rect 47 8 48 12
rect 52 8 53 12
rect 47 7 53 8
rect 55 7 58 13
rect 60 12 66 13
rect 60 8 61 12
rect 65 8 66 12
rect 60 7 66 8
rect 68 7 71 13
rect 73 12 78 13
rect 73 8 74 12
rect 73 7 78 8
rect 88 12 93 14
rect 92 8 93 12
rect 88 7 93 8
rect 95 12 100 14
rect 95 8 96 12
rect 95 7 100 8
<< pdiffusion >>
rect 10 74 11 83
rect 13 74 16 83
rect 18 74 19 83
rect 23 74 24 83
rect 26 74 29 83
rect 31 74 32 83
rect 36 74 37 83
rect 39 74 40 83
rect 44 74 45 83
rect 47 74 48 83
rect 52 74 53 83
rect 55 74 58 83
rect 60 74 61 83
rect 65 74 66 83
rect 68 74 71 83
rect 73 74 74 83
rect 88 82 93 83
rect 92 73 93 82
rect 95 82 100 83
rect 95 73 96 82
<< ndcontact >>
rect 6 8 10 12
rect 19 8 23 12
rect 32 8 36 12
rect 40 8 44 12
rect 48 8 52 12
rect 61 8 65 12
rect 74 8 78 12
rect 88 8 92 12
rect 96 8 100 12
<< pdcontact >>
rect 6 74 10 83
rect 19 74 23 83
rect 32 74 36 83
rect 40 74 44 83
rect 48 74 52 83
rect 61 74 65 83
rect 74 74 78 83
rect 88 73 92 82
rect 96 73 100 82
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
rect 40 -2 44 2
rect 48 -2 52 2
rect 56 -2 60 2
rect 64 -2 68 2
rect 72 -2 76 2
rect 80 -2 84 2
rect 88 -2 92 2
rect 96 -2 100 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
rect 32 88 36 92
rect 40 88 44 92
rect 48 88 52 92
rect 56 88 60 92
rect 64 88 68 92
rect 72 88 76 92
rect 80 88 84 92
rect 88 88 92 92
rect 96 88 100 92
<< polysilicon >>
rect 11 83 13 85
rect 16 83 18 85
rect 24 83 26 85
rect 29 83 31 85
rect 37 83 39 85
rect 45 83 47 85
rect 53 83 55 85
rect 58 83 60 85
rect 66 83 68 85
rect 71 83 73 85
rect 93 83 95 85
rect 11 57 13 74
rect 0 22 2 42
rect 8 30 10 56
rect 16 38 18 74
rect 24 52 26 74
rect 0 20 13 22
rect 11 13 13 20
rect 16 13 18 34
rect 22 50 26 52
rect 22 22 24 50
rect 29 46 31 74
rect 37 53 39 74
rect 45 50 47 74
rect 53 60 55 74
rect 58 73 60 74
rect 58 71 62 73
rect 60 53 62 71
rect 66 59 68 74
rect 71 73 73 74
rect 71 71 78 73
rect 66 57 71 59
rect 60 50 61 53
rect 37 45 39 49
rect 45 48 49 50
rect 37 43 44 45
rect 36 29 38 34
rect 42 29 44 43
rect 47 38 49 48
rect 57 42 58 45
rect 47 35 48 38
rect 56 30 58 42
rect 62 35 64 49
rect 36 27 39 29
rect 42 27 47 29
rect 22 20 26 22
rect 24 13 26 20
rect 29 13 31 26
rect 37 13 39 27
rect 45 13 47 27
rect 53 28 58 30
rect 61 33 64 35
rect 53 13 55 28
rect 61 25 63 33
rect 69 29 71 57
rect 76 46 78 71
rect 84 38 86 56
rect 75 33 76 37
rect 81 36 86 38
rect 58 23 63 25
rect 66 27 71 29
rect 58 13 60 23
rect 66 13 68 27
rect 81 16 83 36
rect 71 14 83 16
rect 93 14 95 73
rect 71 13 73 14
rect 11 5 13 7
rect 16 5 18 7
rect 24 5 26 7
rect 29 5 31 7
rect 37 5 39 7
rect 45 5 47 7
rect 53 5 55 7
rect 58 5 60 7
rect 66 5 68 7
rect 71 5 73 7
rect 93 5 95 7
<< polycontact >>
rect 7 56 11 60
rect 0 42 4 46
rect 14 34 18 38
rect 6 26 10 30
rect 36 49 40 53
rect 51 56 55 60
rect 28 42 32 46
rect 61 49 65 53
rect 24 34 28 38
rect 34 34 38 38
rect 28 26 32 30
rect 53 42 57 46
rect 48 34 52 38
rect 83 56 87 60
rect 75 42 79 46
rect 71 33 75 37
rect 89 27 93 31
<< metal1 >>
rect -2 92 102 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 32 92
rect 36 88 40 92
rect 44 88 48 92
rect 52 88 56 92
rect 60 88 64 92
rect 68 88 72 92
rect 76 88 80 92
rect 84 88 88 92
rect 92 88 96 92
rect 100 88 102 92
rect -2 86 102 88
rect 19 83 23 86
rect 61 83 65 86
rect 6 71 10 74
rect 32 71 36 74
rect 48 71 52 74
rect 74 71 78 74
rect 88 82 92 86
rect 96 82 100 83
rect 6 67 36 71
rect 48 67 78 71
rect 11 56 51 60
rect 55 56 80 60
rect 60 49 61 53
rect 4 42 28 46
rect 32 42 53 46
rect 57 42 75 46
rect 96 41 100 73
rect 38 34 48 38
rect 81 30 89 31
rect 10 26 28 30
rect 44 27 89 30
rect 44 26 85 27
rect 6 16 36 20
rect 6 12 10 16
rect 6 7 10 8
rect 19 12 23 13
rect 19 4 23 8
rect 32 12 36 16
rect 48 16 78 20
rect 32 7 36 8
rect 40 7 44 8
rect 48 12 52 16
rect 48 7 52 8
rect 61 12 65 13
rect 61 4 65 8
rect 74 12 78 16
rect 74 7 78 8
rect 88 12 92 14
rect 88 4 92 8
rect 96 12 100 37
rect 96 7 100 8
rect -2 2 102 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 40 2
rect 44 -2 48 2
rect 52 -2 56 2
rect 60 -2 64 2
rect 68 -2 72 2
rect 76 -2 80 2
rect 84 -2 88 2
rect 92 -2 96 2
rect 100 -2 102 2
rect -2 -4 102 -2
<< m2contact >>
rect 40 74 44 75
rect 40 71 44 74
rect 80 56 83 60
rect 83 56 84 60
rect 32 49 36 53
rect 56 49 60 53
rect 0 42 4 46
rect 16 34 18 38
rect 18 34 20 38
rect 24 34 28 38
rect 48 34 52 38
rect 96 37 100 41
rect 72 33 75 37
rect 75 33 76 37
rect 40 26 44 30
rect 40 12 44 14
rect 40 10 44 12
<< metal2 >>
rect 40 30 44 71
rect 40 14 44 26
rect 40 9 44 10
<< labels >>
rlabel metal1 -1 0 -1 0 3 Gnd!
rlabel m2contact 2 44 2 44 1 s0b
rlabel m2contact 18 36 18 36 1 d0
rlabel m2contact 26 36 26 36 1 d1
rlabel m2contact 34 51 34 51 1 s1
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel m2contact 58 51 58 51 1 d2
rlabel m2contact 82 58 82 58 1 s0
rlabel m2contact 98 39 98 39 1 y
rlabel m2contact 74 35 74 35 1 d3
rlabel m2contact 50 36 50 36 1 s1b
<< end >>
