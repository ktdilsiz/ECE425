magic
tech scmos
timestamp 1484534138
<< nwell >>
rect -6 40 66 96
<< ntransistor >>
rect 8 7 10 13
rect 16 7 18 13
rect 21 7 23 13
rect 29 7 31 13
rect 34 7 36 13
rect 53 7 55 14
<< ptransistor >>
rect 8 74 10 83
rect 16 74 18 83
rect 21 74 23 83
rect 29 74 31 83
rect 34 74 36 83
rect 53 73 55 83
<< ndiffusion >>
rect 3 12 8 13
rect 7 8 8 12
rect 3 7 8 8
rect 10 12 16 13
rect 10 8 11 12
rect 15 8 16 12
rect 10 7 16 8
rect 18 7 21 13
rect 23 7 24 13
rect 28 7 29 13
rect 31 7 34 13
rect 36 12 41 13
rect 36 8 37 12
rect 36 7 41 8
rect 48 12 53 14
rect 52 8 53 12
rect 48 7 53 8
rect 55 12 60 14
rect 55 8 56 12
rect 55 7 60 8
<< pdiffusion >>
rect 7 74 8 83
rect 10 74 11 83
rect 15 74 16 83
rect 18 74 21 83
rect 23 79 24 83
rect 28 79 29 83
rect 23 74 29 79
rect 31 74 34 83
rect 36 74 37 83
rect 48 82 53 83
rect 52 73 53 82
rect 55 82 60 83
rect 55 73 56 82
<< ndcontact >>
rect 3 8 7 12
rect 11 8 15 12
rect 24 7 28 13
rect 37 8 41 12
rect 48 8 52 12
rect 56 8 60 12
<< pdcontact >>
rect 3 74 7 83
rect 11 74 15 83
rect 24 79 28 83
rect 37 74 41 83
rect 48 73 52 82
rect 56 73 60 82
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
rect 40 -2 44 2
rect 48 -2 52 2
rect 56 -2 60 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
rect 32 88 36 92
rect 40 88 44 92
rect 48 88 52 92
rect 56 88 60 92
<< polysilicon >>
rect 8 83 10 85
rect 16 83 18 85
rect 21 83 23 85
rect 29 83 31 85
rect 34 83 36 85
rect 53 83 55 85
rect 8 70 10 74
rect 3 68 10 70
rect 3 55 5 68
rect 16 59 18 74
rect 10 57 18 59
rect 3 16 5 51
rect 10 47 12 57
rect 21 50 23 74
rect 29 73 31 74
rect 18 48 23 50
rect 26 71 31 73
rect 10 22 12 43
rect 18 39 20 48
rect 26 42 28 71
rect 34 62 36 74
rect 34 60 43 62
rect 41 57 43 60
rect 40 53 44 57
rect 24 40 28 42
rect 24 29 26 40
rect 21 27 26 29
rect 29 33 35 35
rect 10 20 18 22
rect 3 14 10 16
rect 8 13 10 14
rect 16 13 18 20
rect 21 13 23 27
rect 29 13 31 33
rect 41 28 43 53
rect 34 26 43 28
rect 34 13 36 26
rect 53 14 55 73
rect 8 5 10 7
rect 16 5 18 7
rect 21 5 23 7
rect 29 5 31 7
rect 34 5 36 7
rect 53 5 55 7
<< polycontact >>
rect 2 51 6 55
rect 9 43 13 47
rect 28 50 32 54
rect 16 35 20 39
rect 32 35 36 39
rect 49 38 53 42
<< metal1 >>
rect -2 92 62 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 32 92
rect 36 88 40 92
rect 44 88 48 92
rect 52 88 56 92
rect 60 88 62 92
rect -2 86 62 88
rect 11 83 15 86
rect 37 83 41 86
rect 24 74 28 79
rect 48 82 52 86
rect 56 82 60 83
rect 6 54 9 55
rect 6 51 28 54
rect 9 50 28 51
rect 28 42 44 46
rect 56 42 60 73
rect 4 35 16 39
rect 20 35 32 39
rect 40 38 49 42
rect 4 12 7 13
rect 3 7 7 8
rect 11 12 15 13
rect 11 4 15 8
rect 37 12 41 13
rect 37 4 41 8
rect 48 12 52 14
rect 48 4 52 8
rect 56 12 60 38
rect 56 7 60 8
rect -2 2 62 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 40 2
rect 44 -2 48 2
rect 52 -2 56 2
rect 60 -2 62 2
rect -2 -4 62 -2
<< m2contact >>
rect 0 74 3 78
rect 3 74 4 78
rect 32 50 36 54
rect 40 53 44 57
rect 8 43 9 47
rect 9 43 12 47
rect 24 42 28 46
rect 0 35 4 39
rect 56 38 60 42
rect 0 12 4 13
rect 0 9 3 12
rect 3 9 4 12
rect 24 9 28 13
<< metal2 >>
rect 0 39 4 74
rect 24 46 28 78
rect 0 13 4 35
rect 24 13 28 42
<< labels >>
rlabel m2contact 10 45 10 45 1 d1
rlabel m2contact 34 52 34 52 1 s
rlabel m2contact 42 55 42 55 1 d0
rlabel m2contact 58 40 58 40 1 y
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel metal1 -1 0 -1 0 2 Gnd!
<< end >>
