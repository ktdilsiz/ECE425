magic
tech scmos
timestamp 1494278851
<< metal1 >>
rect 3961 3850 4007 3851
rect 3965 3846 4007 3850
rect 3961 3845 4007 3846
rect 3968 3550 4006 3551
rect 3972 3546 4006 3550
rect 3968 3544 4006 3546
rect 2904 3275 2960 3276
rect 2904 3271 3965 3275
rect 2904 3267 3961 3271
rect 2904 3262 3965 3267
rect 2904 3261 2960 3262
rect 2904 3212 2916 3261
rect 1105 3200 1208 3207
rect 1105 3176 1109 3200
rect 1119 3080 1124 3200
rect 2205 3198 2916 3212
rect 2920 3237 2935 3239
rect 2920 3235 2941 3237
rect 2920 3230 2935 3235
rect 2940 3230 2941 3235
rect 2920 3228 2941 3230
rect 2920 3185 2935 3228
rect 2176 3173 2935 3185
rect 1104 3074 1124 3080
rect 2920 3030 2935 3173
rect 2929 3021 2935 3030
rect 2945 2998 2960 3261
rect 2964 3235 3972 3237
rect 2964 3230 2965 3235
rect 2970 3231 3968 3235
rect 2970 3230 3972 3231
rect 2964 3228 3972 3230
rect 3815 3134 3965 3135
rect 3815 3130 3961 3134
rect 3815 3127 3965 3130
rect 3815 3043 3972 3045
rect 3815 3039 3968 3043
rect 3815 3037 3972 3039
rect 3815 3003 3965 3005
rect 3815 2999 3961 3003
rect 3815 2997 3965 2999
rect 3815 2913 3972 2915
rect 3815 2909 3968 2913
rect 3815 2907 3972 2909
rect 3815 2873 3965 2875
rect 3815 2869 3961 2873
rect 3815 2867 3965 2869
rect 3815 2783 3972 2785
rect 3815 2779 3968 2783
rect 3815 2777 3972 2779
rect 3815 2743 3965 2745
rect 3815 2739 3961 2743
rect 3815 2737 3965 2739
rect 3815 2654 3972 2655
rect 3815 2650 3968 2654
rect 3815 2647 3972 2650
rect 3910 2484 3965 2486
rect 3910 2480 3961 2484
rect 3910 2478 3965 2480
rect 3958 2394 3972 2396
rect 3958 2390 3968 2394
rect 3958 2388 3972 2390
rect 3910 2375 3965 2376
rect 3910 2371 3961 2375
rect 3910 2368 3965 2371
rect 3958 2284 3972 2286
rect 3958 2280 3968 2284
rect 3958 2278 3972 2280
rect 3910 2264 3965 2266
rect 3910 2260 3961 2264
rect 3910 2258 3965 2260
rect 3958 2174 3972 2176
rect 3958 2170 3968 2174
rect 3958 2168 3972 2170
rect 3910 2155 3965 2156
rect 3910 2151 3961 2155
rect 3910 2148 3965 2151
rect 3958 2064 3972 2066
rect 3958 2060 3968 2064
rect 3958 2058 3972 2060
rect 3910 2044 3965 2046
rect 3910 2040 3961 2044
rect 3910 2038 3965 2040
rect 3958 1954 3972 1956
rect 3958 1950 3968 1954
rect 3958 1948 3972 1950
rect 3910 1934 3965 1936
rect 3910 1930 3961 1934
rect 3910 1928 3965 1930
rect 3958 1844 3972 1846
rect 3958 1840 3968 1844
rect 3958 1838 3972 1840
rect 3910 1824 3965 1826
rect 3910 1820 3961 1824
rect 3910 1818 3965 1820
rect 3958 1734 3972 1736
rect 3958 1730 3968 1734
rect 3958 1728 3972 1730
rect 3910 1715 3965 1716
rect 3910 1711 3961 1715
rect 3910 1708 3965 1711
rect 3958 1624 3972 1626
rect 3958 1620 3968 1624
rect 3958 1618 3972 1620
rect 3910 1604 3965 1606
rect 3910 1600 3961 1604
rect 3910 1598 3965 1600
rect 3958 1514 3972 1516
rect 3958 1510 3968 1514
rect 3958 1508 3972 1510
rect 3910 1494 3965 1496
rect 3910 1490 3961 1494
rect 3910 1488 3965 1490
rect 3958 1404 3972 1406
rect 3958 1400 3968 1404
rect 3958 1398 3972 1400
rect 3910 1384 3965 1386
rect 3910 1380 3961 1384
rect 3910 1378 3965 1380
rect 3958 1294 3972 1296
rect 3958 1290 3968 1294
rect 3958 1288 3972 1290
rect 3910 1274 3965 1276
rect 3910 1270 3961 1274
rect 3910 1268 3965 1270
rect 3958 1184 3972 1186
rect 3958 1180 3968 1184
rect 3958 1178 3972 1180
<< m2contact >>
rect 3961 3846 3965 3850
rect 3968 3546 3972 3550
rect 3961 3267 3965 3271
rect 2935 3230 2940 3235
rect 2920 3021 2929 3030
rect 2965 3230 2970 3235
rect 3968 3231 3972 3235
rect 3961 3130 3965 3134
rect 3968 3039 3972 3043
rect 3961 2999 3965 3003
rect 3968 2909 3972 2913
rect 3961 2869 3965 2873
rect 3968 2779 3972 2783
rect 3961 2739 3965 2743
rect 3968 2650 3972 2654
rect 3961 2480 3965 2484
rect 3968 2390 3972 2394
rect 3961 2371 3965 2375
rect 3968 2280 3972 2284
rect 3961 2260 3965 2264
rect 3968 2170 3972 2174
rect 3961 2151 3965 2155
rect 3968 2060 3972 2064
rect 3961 2040 3965 2044
rect 3968 1950 3972 1954
rect 3961 1930 3965 1934
rect 3968 1840 3972 1844
rect 3961 1820 3965 1824
rect 3968 1730 3972 1734
rect 3961 1711 3965 1715
rect 3968 1620 3972 1624
rect 3961 1600 3965 1604
rect 3968 1510 3972 1514
rect 3961 1490 3965 1494
rect 3968 1400 3972 1404
rect 3961 1380 3965 1384
rect 3968 1290 3972 1294
rect 3961 1270 3965 1274
rect 3968 1180 3972 1184
<< metal2 >>
rect 3961 3850 3965 3962
rect 3961 3271 3965 3846
rect 2933 3235 2990 3238
rect 2933 3230 2935 3235
rect 2940 3230 2965 3235
rect 2970 3230 2990 3235
rect 2933 3228 2990 3230
rect 3961 3134 3965 3267
rect 2920 3030 2935 3032
rect 2929 3021 2935 3030
rect 2920 2992 2935 3021
rect 3961 3003 3965 3130
rect 3961 2873 3965 2999
rect 3961 2743 3965 2869
rect 3961 2484 3965 2739
rect 3961 2375 3965 2480
rect 3961 2264 3965 2371
rect 3961 2155 3965 2260
rect 3961 2044 3965 2151
rect 3961 1934 3965 2040
rect 993 1859 1015 1863
rect 3961 1824 3965 1930
rect 3961 1715 3965 1820
rect 3961 1604 3965 1711
rect 3961 1494 3965 1600
rect 3961 1384 3965 1490
rect 3961 1274 3965 1380
rect 3961 1150 3965 1270
rect 3968 3550 3975 3551
rect 3972 3546 3975 3550
rect 3968 3544 3975 3546
rect 3968 3235 3972 3544
rect 3968 3043 3972 3231
rect 3968 2913 3972 3039
rect 3968 2783 3972 2909
rect 3968 2654 3972 2779
rect 3968 2394 3972 2650
rect 3968 2284 3972 2390
rect 3968 2174 3972 2280
rect 3968 2064 3972 2170
rect 3968 1954 3972 2060
rect 3968 1844 3972 1950
rect 3968 1734 3972 1840
rect 3968 1624 3972 1730
rect 3968 1514 3972 1620
rect 3968 1404 3972 1510
rect 3968 1294 3972 1400
rect 3968 1184 3972 1290
rect 3968 1150 3972 1180
<< m2p >>
rect 1002 1859 1003 1863
use PADFC  PADFC_0
timestamp 949001400
transform 1 0 0 0 1 4000
box 327 -3 1003 673
use PADINC  reset
timestamp 1084294328
transform 1 0 1000 0 1 4000
box -6 -3 303 1000
use PADOUT  adr0
timestamp 1084294529
transform 1 0 1300 0 1 4000
box -6 -3 303 1000
use PADOUT  adr1
timestamp 1084294529
transform 1 0 1600 0 1 4000
box -6 -3 303 1000
use PADOUT  adr2
timestamp 1084294529
transform 1 0 1900 0 1 4000
box -6 -3 303 1000
use PADOUT  adr3
timestamp 1084294529
transform 1 0 2200 0 1 4000
box -6 -3 303 1000
use PADOUT  adr4
timestamp 1084294529
transform 1 0 2500 0 1 4000
box -6 -3 303 1000
use PADOUT  adr5
timestamp 1084294529
transform 1 0 2800 0 1 4000
box -6 -3 303 1000
use PADOUT  adr6
timestamp 1084294529
transform 1 0 3100 0 1 4000
box -6 -3 303 1000
use PADOUT  adr7
timestamp 1084294529
transform 1 0 3400 0 1 4000
box -6 -3 303 1000
use PADOUT  MemWrite
timestamp 1084294529
transform 1 0 3700 0 1 4000
box -6 -3 303 1000
use PADFC  PADFC_3
timestamp 949001400
transform 0 1 4000 -1 0 5000
box 327 -3 1003 673
use PADINC  ph1
timestamp 1084294328
transform 0 -1 1000 1 0 3700
box -6 -3 303 1000
use PADINC  ph2
timestamp 1084294328
transform 0 -1 1000 1 0 3400
box -6 -3 303 1000
use PADVDD  PADVDD_0
timestamp 1084294447
transform 0 1 4000 -1 0 3997
box -3 -3 303 1000
use PADGND  PADGND_0
timestamp 1084294269
transform 0 1 4000 -1 0 3698
box -3 -3 303 1000
use PADINC  memdata7
timestamp 1084294328
transform 0 -1 1000 1 0 3100
box -6 -3 303 1000
use PADINC  memdata6
timestamp 1084294328
transform 0 -1 1000 1 0 2800
box -6 -3 303 1000
use PADINC  memdata5
timestamp 1084294328
transform 0 -1 1000 1 0 2500
box -6 -3 303 1000
use PADINC  memdata4
timestamp 1084294328
transform 0 -1 1000 1 0 2200
box -6 -3 303 1000
use PADINC  memdata3
timestamp 1084294328
transform 0 -1 1000 1 0 1900
box -6 -3 303 1000
use PADINC  memdata2
timestamp 1084294328
transform 0 -1 1000 1 0 1600
box -6 -3 303 1000
use PADOUT  memdata1
timestamp 1084294529
transform 0 -1 1000 1 0 1300
box -6 -3 303 1000
use datapath  datapath_0
timestamp 1494278851
transform 1 0 1219 0 1 1182
box -168 -32 2739 2085
use PADNC  PADNC_9
timestamp 1084294400
transform 0 1 4000 1 0 3100
box -3 -3 303 1000
use PADNC  PADNC_8
timestamp 1084294400
transform 0 1 4000 1 0 2800
box -3 -3 303 1000
use PADNC  PADNC_7
timestamp 1084294400
transform 0 1 4000 1 0 2500
box -3 -3 303 1000
use PADNC  PADNC_6
timestamp 1084294400
transform 0 1 4000 1 0 2200
box -3 -3 303 1000
use PADNC  PADNC_5
timestamp 1084294400
transform 0 1 4000 1 0 1900
box -3 -3 303 1000
use PADNC  PADNC_4
timestamp 1084294400
transform 0 1 4000 1 0 1600
box -3 -3 303 1000
use PADNC  PADNC_3
timestamp 1084294400
transform 0 1 4000 1 0 1300
box -3 -3 303 1000
use PADOUT  memdata0
timestamp 1084294529
transform 0 -1 1000 1 0 1000
box -6 -3 303 1000
use PADFC  PADFC_2
timestamp 949001400
transform 0 -1 1000 1 0 0
box 327 -3 1003 673
use PADOUT  writedata0
timestamp 1084294529
transform -1 0 1300 0 -1 1000
box -6 -3 303 1000
use PADOUT  writedata1
timestamp 1084294529
transform -1 0 1600 0 -1 1000
box -6 -3 303 1000
use PADOUT  writedata2
timestamp 1084294529
transform -1 0 1900 0 -1 1000
box -6 -3 303 1000
use PADOUT  writedata3
timestamp 1084294529
transform -1 0 2200 0 -1 1000
box -6 -3 303 1000
use PADOUT  writedata4
timestamp 1084294529
transform -1 0 2500 0 -1 1000
box -6 -3 303 1000
use PADOUT  writedata5
timestamp 1084294529
transform -1 0 2800 0 -1 1000
box -6 -3 303 1000
use PADOUT  writedata6
timestamp 1084294529
transform -1 0 3100 0 -1 1000
box -6 -3 303 1000
use PADOUT  writedata7
timestamp 1084294529
transform -1 0 3400 0 -1 1000
box -6 -3 303 1000
use PADNC  PADNC_0
timestamp 1084294400
transform 1 0 3400 0 -1 1000
box -3 -3 303 1000
use PADNC  PADNC_1
timestamp 1084294400
transform 0 1 4000 1 0 1000
box -3 -3 303 1000
use PADFC  PADFC_1
timestamp 949001400
transform -1 0 4998 0 -1 1000
box 327 -3 1003 673
use PADNC  PADNC_2
timestamp 1084294400
transform 1 0 3700 0 -1 1000
box -3 -3 303 1000
<< end >>
