magic
tech scmos
timestamp 1494266977
<< nwell >>
rect -8 48 32 105
<< ntransistor >>
rect 7 6 9 16
rect 15 6 17 16
<< ptransistor >>
rect 7 54 9 94
rect 12 54 14 94
<< ndiffusion >>
rect 2 15 7 16
rect 6 6 7 15
rect 9 15 15 16
rect 9 6 10 15
rect 14 6 15 15
rect 17 15 22 16
rect 17 6 18 15
<< pdiffusion >>
rect 2 93 7 94
rect 6 54 7 93
rect 9 54 12 94
rect 14 93 19 94
rect 14 54 15 93
<< ndcontact >>
rect 2 6 6 15
rect 10 6 14 15
rect 18 6 22 15
<< pdcontact >>
rect 2 54 6 93
rect 15 54 19 93
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 12 94 14 96
rect 7 23 9 54
rect 12 53 14 54
rect 12 51 17 53
rect 6 19 9 23
rect 7 16 9 19
rect 15 47 18 51
rect 15 16 17 47
rect 7 4 9 6
rect 15 4 17 6
<< polycontact >>
rect 2 19 6 23
rect 18 47 22 51
<< metal1 >>
rect -2 102 26 103
rect 2 98 14 102
rect 18 98 26 102
rect -2 97 26 98
rect 2 93 6 97
rect 15 93 19 94
rect 10 54 15 58
rect 11 37 14 54
rect 18 43 22 47
rect 10 33 14 37
rect 2 23 6 27
rect 11 16 14 33
rect 2 15 6 16
rect 10 15 14 16
rect 18 15 22 16
rect 2 3 6 6
rect 18 3 22 6
rect -2 2 26 3
rect 2 -2 14 2
rect 18 -2 26 2
rect -2 -3 26 -2
<< labels >>
flabel metal1 4 100 4 100 4 FreeSans 26 0 0 0 vdd
flabel metal1 20 45 20 45 4 FreeSans 26 0 0 0 B
flabel metal1 4 0 4 0 4 FreeSans 26 0 0 0 gnd
flabel metal1 12 35 12 35 4 FreeSans 26 0 0 0 Y
flabel metal1 4 25 4 25 4 FreeSans 26 0 0 0 A
<< end >>
