magic
tech scmos
timestamp 1484419682
<< nwell >>
rect -6 40 34 96
<< ntransistor >>
rect 5 7 7 14
rect 13 7 15 13
rect 21 7 23 13
<< ptransistor >>
rect 5 73 7 83
rect 13 71 15 83
rect 18 71 20 83
<< ndiffusion >>
rect 0 12 5 14
rect 4 8 5 12
rect 0 7 5 8
rect 7 13 12 14
rect 7 12 13 13
rect 7 8 8 12
rect 12 8 13 12
rect 7 7 13 8
rect 15 12 21 13
rect 15 8 16 12
rect 20 8 21 12
rect 15 7 21 8
rect 23 12 28 13
rect 23 8 24 12
rect 23 7 28 8
<< pdiffusion >>
rect 0 82 5 83
rect 4 73 5 82
rect 7 82 13 83
rect 7 73 8 82
rect 12 73 13 82
rect 10 71 13 73
rect 15 71 18 83
rect 20 81 25 83
rect 20 72 21 81
rect 20 71 25 72
<< ndcontact >>
rect 0 8 4 12
rect 8 8 12 12
rect 16 8 20 12
rect 24 8 28 12
<< pdcontact >>
rect 0 73 4 82
rect 8 73 12 82
rect 21 72 25 81
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
<< polysilicon >>
rect 5 83 7 85
rect 13 83 15 85
rect 18 83 20 85
rect 5 41 7 73
rect 13 48 15 71
rect 18 57 20 71
rect 18 55 28 57
rect 5 39 11 41
rect 5 14 7 39
rect 19 34 21 50
rect 13 32 21 34
rect 13 13 15 32
rect 26 26 28 55
rect 25 16 28 22
rect 21 14 28 16
rect 21 13 23 14
rect 5 5 7 7
rect 13 5 15 7
rect 21 5 23 7
<< polycontact >>
rect 15 47 19 51
rect 11 38 15 42
rect 24 22 28 26
<< metal1 >>
rect -2 92 30 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 30 92
rect -2 86 30 88
rect 0 82 4 83
rect 8 82 12 86
rect 21 81 25 83
rect 0 42 4 73
rect 21 59 25 72
rect 21 55 28 59
rect 24 42 28 55
rect 15 38 28 42
rect 0 12 4 38
rect 0 7 4 8
rect 8 12 12 14
rect 8 4 12 8
rect 16 12 20 38
rect 16 7 20 8
rect 24 12 28 13
rect 24 4 28 8
rect -2 2 30 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 30 2
rect -2 -4 30 -2
<< m2contact >>
rect 17 47 19 51
rect 19 47 21 51
rect 0 38 4 42
rect 24 22 28 26
<< metal2 >>
rect 16 47 17 51
<< labels >>
rlabel m2contact 19 49 19 49 1 a
rlabel m2contact 26 24 26 24 1 b
rlabel m2contact 2 40 2 40 1 y
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel metal1 -1 0 -1 0 3 Gnd!
<< end >>
