magic
tech scmos
timestamp 1487713933
<< nwell >>
rect -6 40 50 96
<< ntransistor >>
rect 5 24 7 30
rect 10 24 12 30
rect 18 24 20 30
rect 23 24 25 30
rect 31 23 33 30
<< ptransistor >>
rect 29 76 39 78
rect 5 54 7 63
rect 13 54 15 63
rect 21 54 23 63
rect 29 54 31 63
<< ndiffusion >>
rect 0 29 5 30
rect 4 25 5 29
rect 0 24 5 25
rect 7 24 10 30
rect 12 29 18 30
rect 12 25 13 29
rect 17 25 18 29
rect 12 24 18 25
rect 20 24 23 30
rect 25 28 31 30
rect 25 24 26 28
rect 30 24 31 28
rect 26 23 31 24
rect 33 28 38 30
rect 33 24 34 28
rect 33 23 38 24
<< pdiffusion >>
rect 38 79 39 83
rect 29 78 39 79
rect 29 75 39 76
rect 38 71 39 75
rect 4 54 5 63
rect 7 54 8 63
rect 12 54 13 63
rect 15 54 16 63
rect 20 54 21 63
rect 23 59 29 63
rect 23 55 24 59
rect 28 55 29 59
rect 23 54 29 55
rect 31 54 32 63
<< ndcontact >>
rect 0 25 4 29
rect 13 25 17 29
rect 26 24 30 28
rect 34 24 38 28
<< pdcontact >>
rect 29 79 38 83
rect 29 71 38 75
rect 0 54 4 63
rect 8 54 12 63
rect 16 54 20 63
rect 24 55 28 59
rect 32 54 36 63
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
rect 40 -2 44 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
rect 32 88 36 92
rect 40 88 44 92
<< polysilicon >>
rect 27 76 29 78
rect 39 76 42 78
rect 5 63 7 65
rect 13 63 15 65
rect 21 63 23 65
rect 29 63 31 65
rect 5 53 7 54
rect 13 53 15 54
rect 21 53 23 54
rect 2 51 7 53
rect 10 51 15 53
rect 18 51 23 53
rect 29 53 31 54
rect 29 51 34 53
rect 2 44 4 51
rect 10 44 12 51
rect 18 44 20 51
rect 32 48 34 51
rect 2 33 4 40
rect 2 31 7 33
rect 5 30 7 31
rect 10 30 12 40
rect 18 30 20 40
rect 26 45 32 47
rect 26 35 28 45
rect 23 33 28 35
rect 31 33 32 35
rect 40 36 42 76
rect 36 34 42 36
rect 23 30 25 33
rect 31 30 33 33
rect 5 22 7 24
rect 10 22 12 24
rect 18 22 20 24
rect 23 22 25 24
rect 31 21 33 23
<< polycontact >>
rect 0 40 4 44
rect 8 40 12 44
rect 16 40 20 44
rect 32 44 36 48
rect 32 33 36 37
<< metal1 >>
rect -2 92 46 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 32 92
rect 36 88 40 92
rect 44 88 46 92
rect -2 86 46 88
rect 8 63 12 86
rect 35 83 39 86
rect 38 79 39 83
rect 38 71 44 75
rect 16 64 36 68
rect 16 63 20 64
rect 32 63 36 64
rect 0 51 4 54
rect 16 51 20 54
rect 0 47 20 51
rect 24 59 28 61
rect 24 37 28 55
rect 40 44 44 71
rect 13 33 32 37
rect 0 29 4 30
rect 0 4 4 25
rect 13 29 17 33
rect 40 30 44 40
rect 13 24 17 25
rect 26 28 30 30
rect 26 4 30 24
rect 34 28 44 30
rect 38 26 44 28
rect 34 23 38 24
rect -2 2 46 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 40 2
rect 44 -2 46 2
rect -2 -4 46 -2
<< m2contact >>
rect 0 40 4 44
rect 8 40 12 44
rect 16 40 20 44
rect 32 44 36 48
rect 40 40 44 44
<< labels >>
rlabel metal1 -1 0 -1 0 3 Gnd!
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel m2contact 42 42 42 42 1 y
rlabel m2contact 2 42 2 42 1 a
rlabel m2contact 10 42 10 42 1 b
rlabel m2contact 18 42 18 42 1 c
rlabel m2contact 34 46 34 46 1 d
<< end >>
