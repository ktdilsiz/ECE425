magic
tech scmos
timestamp 1484514831
<< nwell >>
rect -6 40 82 96
<< ntransistor >>
rect 5 7 7 13
rect 10 7 12 13
rect 18 7 20 13
rect 23 7 25 13
rect 31 7 33 13
rect 39 7 41 13
rect 44 7 46 13
rect 62 12 69 14
<< ptransistor >>
rect 5 74 7 83
rect 10 74 12 83
rect 18 74 20 83
rect 23 74 25 83
rect 31 74 33 83
rect 39 74 41 83
rect 44 74 46 83
rect 59 73 69 75
<< ndiffusion >>
rect 62 15 63 19
rect 67 15 69 19
rect 62 14 69 15
rect 0 12 5 13
rect 4 8 5 12
rect 0 7 5 8
rect 7 7 10 13
rect 12 12 18 13
rect 12 8 13 12
rect 17 8 18 12
rect 12 7 18 8
rect 20 7 23 13
rect 25 12 31 13
rect 25 8 26 12
rect 30 8 31 12
rect 25 7 31 8
rect 33 12 39 13
rect 33 8 34 12
rect 38 8 39 12
rect 33 7 39 8
rect 41 7 44 13
rect 46 12 51 13
rect 46 8 47 12
rect 46 7 51 8
rect 62 11 69 12
rect 62 7 63 11
rect 67 7 69 11
<< pdiffusion >>
rect 4 74 5 83
rect 7 74 10 83
rect 12 74 13 83
rect 17 74 18 83
rect 20 74 23 83
rect 25 74 26 83
rect 30 74 31 83
rect 33 74 34 83
rect 38 74 39 83
rect 41 74 44 83
rect 46 74 47 83
rect 68 76 69 80
rect 59 75 69 76
rect 59 72 69 73
rect 68 68 69 72
<< ndcontact >>
rect 63 15 67 19
rect 0 8 4 12
rect 13 8 17 12
rect 26 8 30 12
rect 34 8 38 12
rect 47 8 51 12
rect 63 7 67 11
<< pdcontact >>
rect 0 74 4 83
rect 13 74 17 83
rect 26 74 30 83
rect 34 74 38 83
rect 47 74 51 83
rect 59 76 68 80
rect 59 68 68 72
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
rect 40 -2 44 2
rect 48 -2 52 2
rect 56 -2 60 2
rect 64 -2 68 2
rect 72 -2 76 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
rect 32 88 36 92
rect 40 88 44 92
rect 48 88 52 92
rect 56 88 60 92
rect 64 88 68 92
rect 72 88 76 92
<< polysilicon >>
rect 5 83 7 85
rect 10 83 12 85
rect 18 83 20 85
rect 23 83 25 85
rect 31 83 33 85
rect 39 83 41 85
rect 44 83 46 85
rect 5 64 7 74
rect 0 62 7 64
rect 0 52 2 62
rect 10 58 12 74
rect 18 64 20 74
rect 9 56 12 58
rect 16 62 20 64
rect 0 26 2 48
rect 9 43 11 56
rect 16 52 18 62
rect 23 59 25 74
rect 31 73 33 74
rect 31 71 36 73
rect 23 57 30 59
rect 28 49 30 57
rect 34 54 36 71
rect 39 59 41 74
rect 44 64 46 74
rect 57 73 59 75
rect 69 73 72 75
rect 44 62 59 64
rect 70 62 72 73
rect 39 57 50 59
rect 34 52 42 54
rect 16 32 18 48
rect 28 47 35 49
rect 23 32 25 39
rect 33 35 35 47
rect 40 43 42 52
rect 48 52 50 57
rect 57 52 59 62
rect 67 58 72 62
rect 60 48 65 51
rect 13 30 18 32
rect 21 30 25 32
rect 29 33 35 35
rect 48 34 50 48
rect 0 24 7 26
rect 5 13 7 24
rect 13 16 15 30
rect 21 27 23 30
rect 29 27 31 33
rect 44 32 50 34
rect 44 30 46 32
rect 10 14 15 16
rect 18 25 23 27
rect 26 25 31 27
rect 34 28 46 30
rect 55 28 57 39
rect 10 13 12 14
rect 18 13 20 25
rect 26 16 28 25
rect 34 22 36 28
rect 53 26 57 28
rect 53 25 55 26
rect 23 14 28 16
rect 31 20 36 22
rect 39 23 55 25
rect 23 13 25 14
rect 31 13 33 20
rect 39 13 41 23
rect 63 22 65 48
rect 59 20 65 22
rect 44 18 61 20
rect 44 13 46 18
rect 70 14 72 58
rect 60 12 62 14
rect 69 12 72 14
rect 5 5 7 7
rect 10 5 12 7
rect 18 5 20 7
rect 23 5 25 7
rect 31 5 33 7
rect 39 5 41 7
rect 44 5 46 7
<< polycontact >>
rect 0 48 4 52
rect 16 48 20 52
rect 24 48 28 52
rect 8 39 12 43
rect 22 39 26 43
rect 63 58 67 62
rect 48 48 52 52
rect 56 48 60 52
rect 40 39 44 43
rect 54 39 58 43
<< metal1 >>
rect -2 92 78 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 32 92
rect 36 88 40 92
rect 44 88 48 92
rect 52 88 56 92
rect 60 88 64 92
rect 68 88 72 92
rect 76 88 78 92
rect -2 86 78 88
rect 13 83 17 86
rect 47 83 51 86
rect 0 70 4 74
rect 26 70 30 74
rect 0 66 30 70
rect 62 80 66 86
rect 68 76 69 80
rect 0 58 4 66
rect 34 62 38 74
rect 68 68 76 72
rect 34 58 63 62
rect 12 39 22 43
rect 44 39 54 43
rect 63 28 67 58
rect 34 24 67 28
rect 72 42 76 68
rect 0 17 30 21
rect 0 12 4 17
rect 0 7 4 8
rect 13 12 17 13
rect 13 4 17 8
rect 26 12 30 17
rect 26 7 30 8
rect 34 12 38 24
rect 72 19 76 38
rect 62 15 63 19
rect 67 15 76 19
rect 34 7 38 8
rect 47 12 51 13
rect 47 4 51 8
rect 62 7 63 11
rect 67 7 69 11
rect 63 4 67 7
rect -2 2 78 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 40 2
rect 44 -2 48 2
rect 52 -2 56 2
rect 60 -2 64 2
rect 68 -2 72 2
rect 76 -2 78 2
rect -2 -4 78 -2
<< m2contact >>
rect 0 48 4 52
rect 16 48 20 52
rect 24 48 28 52
rect 48 48 52 52
rect 56 48 60 52
rect 8 39 12 43
rect 40 39 44 43
rect 72 38 76 42
<< labels >>
rlabel m2contact 2 50 2 50 1 s0
rlabel m2contact 18 50 18 50 1 d1
rlabel m2contact 26 50 26 50 1 s0b
rlabel m2contact 50 50 50 50 1 s1b
rlabel m2contact 58 50 58 50 1 d2
rlabel m2contact 74 40 74 40 1 y
rlabel m2contact 42 41 42 41 1 s1
rlabel m2contact 10 41 10 41 1 d0
rlabel metal1 -1 89 -1 89 3 Vdd!
rlabel metal1 -1 0 -1 0 2 Gnd!
<< end >>
