magic
tech scmos
timestamp 1487715319
<< nwell >>
rect -4 40 44 96
<< ntransistor >>
rect 7 7 9 28
rect 12 7 14 28
rect 20 7 22 21
<< ptransistor >>
rect 7 46 9 83
rect 15 46 17 83
rect 23 46 25 83
<< ndiffusion >>
rect 2 27 7 28
rect 6 8 7 27
rect 2 7 7 8
rect 9 7 12 28
rect 14 27 19 28
rect 14 8 15 27
rect 19 8 20 21
rect 14 7 20 8
rect 22 7 23 21
<< pdiffusion >>
rect 2 81 7 83
rect 6 47 7 81
rect 2 46 7 47
rect 9 82 15 83
rect 9 48 10 82
rect 14 48 15 82
rect 9 46 15 48
rect 17 81 23 83
rect 17 47 18 81
rect 22 47 23 81
rect 17 46 23 47
rect 25 81 30 83
rect 25 47 26 81
rect 25 46 30 47
<< ndcontact >>
rect 2 8 6 27
rect 15 8 19 27
rect 23 7 27 21
<< pdcontact >>
rect 2 47 6 81
rect 10 48 14 82
rect 18 47 22 81
rect 26 47 30 81
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 88 6 92
rect 10 88 14 92
rect 18 88 22 92
rect 26 88 30 92
rect 34 88 38 92
<< polysilicon >>
rect 7 83 9 85
rect 15 83 17 85
rect 23 83 25 85
rect 7 45 9 46
rect 2 43 9 45
rect 2 36 4 43
rect 15 36 17 46
rect 23 45 25 46
rect 23 43 26 45
rect 2 30 9 32
rect 7 28 9 30
rect 12 30 17 32
rect 24 36 26 43
rect 34 32 38 36
rect 12 28 14 30
rect 24 24 26 32
rect 20 22 26 24
rect 20 21 22 22
rect 7 5 9 7
rect 12 5 14 7
rect 20 5 22 7
<< polycontact >>
rect 2 32 6 36
rect 13 32 17 36
rect 24 32 28 36
<< metal1 >>
rect 0 92 40 94
rect 0 88 2 92
rect 6 88 10 92
rect 14 88 18 92
rect 22 88 26 92
rect 30 88 34 92
rect 38 88 40 92
rect 0 86 40 88
rect 2 81 6 83
rect 10 82 14 86
rect 10 47 14 48
rect 18 81 22 83
rect 2 44 6 47
rect 18 44 22 47
rect 2 40 22 44
rect 26 81 30 83
rect 26 44 30 47
rect 26 40 38 44
rect 34 36 38 40
rect 34 28 38 32
rect 2 27 6 28
rect 2 4 6 8
rect 15 27 38 28
rect 19 24 38 27
rect 15 7 19 8
rect 23 4 27 7
rect 0 2 40 4
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -4 40 -2
<< m2contact >>
rect 2 32 6 36
rect 10 32 13 36
rect 13 32 14 36
rect 26 32 28 36
rect 28 32 30 36
rect 34 32 38 36
<< labels >>
rlabel metal1 1 0 1 0 2 Gnd!
rlabel metal1 1 90 1 90 3 Vdd!
rlabel m2contact 4 34 4 34 1 a
rlabel m2contact 12 34 12 34 1 b
rlabel m2contact 28 34 28 34 1 c
rlabel m2contact 36 34 36 34 1 y
<< end >>
