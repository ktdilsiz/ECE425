magic
tech scmos
timestamp 1486493186
<< nwell >>
rect -6 40 34 96
<< ntransistor >>
rect 5 9 7 25
rect 10 9 12 25
rect 15 9 17 25
<< ptransistor >>
rect 5 70 7 83
rect 13 70 15 83
rect 21 70 23 83
<< ndiffusion >>
rect 4 9 5 25
rect 7 9 10 25
rect 12 9 15 25
rect 17 9 18 25
<< pdiffusion >>
rect 4 70 5 83
rect 7 70 8 83
rect 12 70 13 83
rect 15 70 16 83
rect 20 70 21 83
rect 23 70 24 83
<< ndcontact >>
rect 0 9 4 25
rect 18 9 22 25
<< pdcontact >>
rect 0 70 4 83
rect 8 70 12 83
rect 16 70 20 83
rect 24 70 28 83
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
<< polysilicon >>
rect 5 83 7 85
rect 13 83 15 85
rect 21 83 23 85
rect 5 67 7 70
rect 13 69 15 70
rect 1 65 7 67
rect 10 67 15 69
rect 1 47 3 65
rect 10 47 12 67
rect 21 60 23 70
rect 20 58 23 60
rect 1 31 3 43
rect 1 29 7 31
rect 5 25 7 29
rect 10 25 12 43
rect 20 31 22 58
rect 15 29 22 31
rect 15 25 17 29
rect 5 7 7 9
rect 10 7 12 9
rect 15 7 17 9
<< polycontact >>
rect 0 43 4 47
rect 8 43 12 47
rect 16 43 20 47
<< metal1 >>
rect -2 92 30 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 30 92
rect -2 86 30 88
rect 0 83 4 86
rect 0 69 4 70
rect 8 66 12 70
rect 24 66 28 70
rect 8 62 28 66
rect 24 47 28 62
rect 24 27 28 43
rect 0 25 4 27
rect 0 4 4 9
rect 18 25 28 27
rect 22 23 28 25
rect 18 7 22 9
rect -2 2 30 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 30 2
rect -2 -4 30 -2
<< m2contact >>
rect 0 43 4 47
rect 8 43 12 47
rect 16 43 20 47
rect 24 43 28 47
<< labels >>
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel metal1 -1 0 -1 0 2 Gnd!
rlabel m2contact 2 45 2 45 1 A
rlabel m2contact 10 45 10 45 1 B
rlabel m2contact 18 45 18 45 1 C
rlabel m2contact 26 45 26 45 1 Y
<< end >>
