magic
tech scmos
timestamp 1492544733
<< metal1 >>
rect -350 151 -12 155
rect -8 151 253 155
rect 257 151 258 155
rect -350 144 -60 148
rect -56 144 221 148
rect 225 144 258 148
rect -350 137 -108 141
rect -104 137 189 141
rect 193 137 258 141
rect -350 130 -156 134
rect -152 130 157 134
rect 161 130 258 134
rect -350 123 -204 127
rect -200 123 125 127
rect 129 123 258 127
rect -350 116 -252 120
rect -248 116 93 120
rect 97 116 258 120
rect -350 109 -300 113
rect -296 109 61 113
rect 65 109 258 113
rect -350 102 -348 106
rect -344 102 -261 106
rect -257 102 20 106
rect 24 102 258 106
<< m2contact >>
rect -12 151 -8 155
rect 253 151 257 155
rect -60 144 -56 148
rect 221 144 225 148
rect -108 137 -104 141
rect 189 137 193 141
rect -156 130 -152 134
rect 157 130 161 134
rect -204 123 -200 127
rect 125 123 129 127
rect -252 116 -248 120
rect 93 116 97 120
rect -300 109 -296 113
rect 61 109 65 113
rect -348 102 -344 106
rect -261 102 -257 106
rect 20 102 24 106
rect -316 -89 -312 -85
rect -308 -89 -304 -85
rect -330 -97 -326 -93
<< metal2 >>
rect -348 49 -344 102
rect -324 -16 -320 62
rect -316 -7 -312 51
rect -300 49 -296 109
rect -316 -85 -312 -20
rect -308 -85 -304 -29
rect -300 -89 -296 -11
rect -276 -16 -272 62
rect -268 -7 -264 51
rect -261 -62 -257 102
rect -252 49 -248 116
rect -228 -16 -224 62
rect -220 -7 -216 51
rect -204 49 -200 123
rect -180 -16 -176 62
rect -172 -7 -168 51
rect -156 49 -152 130
rect -132 -16 -128 62
rect -124 -7 -120 51
rect -108 49 -104 137
rect -84 -16 -80 62
rect -76 -7 -72 51
rect -60 49 -56 144
rect -36 -16 -32 62
rect -28 -7 -24 51
rect -12 49 -8 151
rect 12 -16 16 62
rect 20 47 24 102
rect 61 64 65 109
rect 93 64 97 116
rect 125 64 129 123
rect 157 64 161 130
rect 189 64 193 137
rect 221 64 225 144
rect 253 64 257 151
rect 52 -16 56 37
rect 84 -16 88 37
rect 116 -16 120 37
rect 148 -16 152 37
rect 180 -16 184 37
rect 212 -16 216 37
rect 244 -16 248 37
rect -124 -211 -120 -90
rect -92 -213 -88 -90
rect -76 -211 -72 -90
rect -44 -213 -40 -90
rect -28 -211 -24 -90
rect 4 -213 8 -90
rect 20 -211 24 -90
rect 52 -213 56 -90
rect 68 -211 72 -90
rect 100 -213 104 -90
rect 116 -211 120 -90
rect 148 -213 152 -90
rect 164 -211 168 -90
rect 196 -213 200 -90
rect 212 -211 216 -90
rect 244 -213 248 -90
rect -84 -216 -80 -215
rect -124 -341 -120 -220
rect -92 -343 -88 -220
rect -76 -341 -72 -220
rect -44 -343 -40 -220
rect -28 -341 -24 -220
rect 4 -343 8 -220
rect 20 -341 24 -220
rect 52 -343 56 -220
rect 68 -341 72 -220
rect 100 -343 104 -220
rect 116 -341 120 -220
rect 148 -343 152 -220
rect 164 -341 168 -220
rect 196 -343 200 -220
rect 212 -341 216 -220
rect 244 -343 248 -220
<< m3contact >>
rect -316 -11 -312 -7
rect -300 -11 -296 -7
rect -324 -20 -320 -16
rect -316 -20 -312 -16
rect -308 -29 -304 -25
rect -268 -11 -264 -7
rect -276 -20 -272 -16
rect -220 -11 -216 -7
rect -228 -20 -224 -16
rect -172 -11 -168 -7
rect -180 -20 -176 -16
rect -124 -11 -120 -7
rect -132 -20 -128 -16
rect -76 -11 -72 -7
rect -84 -20 -80 -16
rect -28 -11 -24 -7
rect -36 -20 -32 -16
rect 12 -20 16 -16
rect 52 -20 56 -16
rect 84 -20 88 -16
rect 116 -20 120 -16
rect 148 -20 152 -16
rect 180 -20 184 -16
rect 212 -20 216 -16
rect 244 -20 248 -16
rect -261 -66 -257 -62
rect -132 -90 -128 -86
rect -124 -90 -120 -86
rect -330 -97 -326 -93
rect -284 -97 -280 -93
rect -92 -90 -88 -86
rect -84 -90 -80 -86
rect -76 -90 -72 -86
rect -44 -90 -40 -86
rect -36 -90 -32 -86
rect -28 -90 -24 -86
rect 4 -90 8 -86
rect 12 -90 16 -86
rect 20 -90 24 -86
rect 52 -90 56 -86
rect 60 -90 64 -86
rect 68 -90 72 -86
rect 100 -90 104 -86
rect 108 -90 112 -86
rect 116 -90 120 -86
rect 148 -90 152 -86
rect 156 -90 160 -86
rect 164 -90 168 -86
rect 196 -90 200 -86
rect 204 -90 208 -86
rect 212 -90 216 -86
rect 244 -90 248 -86
rect -132 -220 -128 -216
rect -124 -220 -120 -216
rect -92 -220 -88 -216
rect -84 -220 -80 -216
rect -76 -220 -72 -216
rect -44 -220 -40 -216
rect -36 -220 -32 -216
rect -28 -220 -24 -216
rect 4 -220 8 -216
rect 12 -220 16 -216
rect 20 -220 24 -216
rect 52 -220 56 -216
rect 60 -220 64 -216
rect 68 -220 72 -216
rect 100 -220 104 -216
rect 108 -220 112 -216
rect 116 -220 120 -216
rect 148 -220 152 -216
rect 156 -220 160 -216
rect 164 -220 168 -216
rect 196 -220 200 -216
rect 204 -220 208 -216
rect 212 -220 216 -216
rect 244 -220 248 -216
<< metal3 >>
rect -348 -7 20 -6
rect -348 -11 -316 -7
rect -312 -11 -300 -7
rect -296 -11 -268 -7
rect -264 -11 -220 -7
rect -216 -11 -172 -7
rect -168 -11 -124 -7
rect -120 -11 -76 -7
rect -72 -11 -28 -7
rect -24 -11 20 -7
rect -348 -12 20 -11
rect -325 -16 256 -15
rect -325 -20 -324 -16
rect -320 -20 -316 -16
rect -312 -20 -276 -16
rect -272 -20 -228 -16
rect -224 -20 -180 -16
rect -176 -20 -132 -16
rect -128 -20 -84 -16
rect -80 -20 -36 -16
rect -32 -20 12 -16
rect 16 -20 52 -16
rect 56 -20 84 -16
rect 88 -20 116 -16
rect 120 -20 148 -16
rect 152 -20 180 -16
rect 184 -20 212 -16
rect 216 -20 244 -16
rect 248 -20 256 -16
rect -325 -21 256 -20
rect -322 -25 -293 -24
rect -322 -29 -308 -25
rect -304 -29 -293 -25
rect -322 -30 -293 -29
rect -276 -62 -256 -61
rect -276 -66 -261 -62
rect -257 -66 -256 -62
rect -276 -67 -256 -66
rect -133 -86 -119 -85
rect -133 -90 -132 -86
rect -128 -90 -124 -86
rect -120 -90 -119 -86
rect -133 -91 -119 -90
rect -93 -86 -71 -85
rect -93 -90 -92 -86
rect -88 -90 -84 -86
rect -80 -90 -76 -86
rect -72 -90 -71 -86
rect -93 -91 -71 -90
rect -45 -86 -23 -85
rect -45 -90 -44 -86
rect -40 -90 -36 -86
rect -32 -90 -28 -86
rect -24 -90 -23 -86
rect -45 -91 -23 -90
rect 3 -86 25 -85
rect 3 -90 4 -86
rect 8 -90 12 -86
rect 16 -90 20 -86
rect 24 -90 25 -86
rect 3 -91 25 -90
rect 51 -86 73 -85
rect 51 -90 52 -86
rect 56 -90 60 -86
rect 64 -90 68 -86
rect 72 -90 73 -86
rect 51 -91 73 -90
rect 99 -86 121 -85
rect 99 -90 100 -86
rect 104 -90 108 -86
rect 112 -90 116 -86
rect 120 -90 121 -86
rect 99 -91 121 -90
rect 147 -86 169 -85
rect 147 -90 148 -86
rect 152 -90 156 -86
rect 160 -90 164 -86
rect 168 -90 169 -86
rect 147 -91 169 -90
rect 195 -86 217 -85
rect 195 -90 196 -86
rect 200 -90 204 -86
rect 208 -90 212 -86
rect 216 -90 217 -86
rect 195 -91 217 -90
rect 243 -86 251 -85
rect 243 -90 244 -86
rect 248 -90 251 -86
rect 243 -91 251 -90
rect -331 -93 -279 -92
rect -331 -97 -330 -93
rect -326 -97 -284 -93
rect -280 -97 -279 -93
rect -331 -98 -279 -97
rect -133 -216 -119 -215
rect -133 -220 -132 -216
rect -128 -220 -124 -216
rect -120 -220 -119 -216
rect -133 -221 -119 -220
rect -93 -216 -71 -215
rect -93 -220 -92 -216
rect -88 -220 -84 -216
rect -80 -220 -76 -216
rect -72 -220 -71 -216
rect -93 -221 -71 -220
rect -45 -216 -23 -215
rect -45 -220 -44 -216
rect -40 -220 -36 -216
rect -32 -220 -28 -216
rect -24 -220 -23 -216
rect -45 -221 -23 -220
rect 3 -216 25 -215
rect 3 -220 4 -216
rect 8 -220 12 -216
rect 16 -220 20 -216
rect 24 -220 25 -216
rect 3 -221 25 -220
rect 51 -216 73 -215
rect 51 -220 52 -216
rect 56 -220 60 -216
rect 64 -220 68 -216
rect 72 -220 73 -216
rect 51 -221 73 -220
rect 99 -216 121 -215
rect 99 -220 100 -216
rect 104 -220 108 -216
rect 112 -220 116 -216
rect 120 -220 121 -216
rect 99 -221 121 -220
rect 147 -216 169 -215
rect 147 -220 148 -216
rect 152 -220 156 -216
rect 160 -220 164 -216
rect 168 -220 169 -216
rect 147 -221 169 -220
rect 195 -216 217 -215
rect 195 -220 196 -216
rect 200 -220 204 -216
rect 208 -220 212 -216
rect 216 -220 217 -216
rect 195 -221 217 -220
rect 243 -216 251 -215
rect 243 -220 244 -216
rect 248 -220 251 -216
rect 243 -221 251 -220
use mux2_dp_1x  mux2_dp_1x_0
timestamp 1484435125
transform 1 0 -348 0 1 3
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_1
timestamp 1484435125
transform 1 0 -300 0 1 3
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_2
timestamp 1484435125
transform 1 0 -252 0 1 3
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_3
timestamp 1484435125
transform 1 0 -204 0 1 3
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_4
timestamp 1484435125
transform 1 0 -156 0 1 3
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_5
timestamp 1484435125
transform 1 0 -108 0 1 3
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_6
timestamp 1484435125
transform 1 0 -60 0 1 3
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_7
timestamp 1484435125
transform 1 0 -12 0 1 3
box -6 -4 50 96
use and2_1x  and2_1x_0
timestamp 1484419738
transform 1 0 36 0 1 3
box -6 -4 34 96
use and2_1x  and2_1x_1
timestamp 1484419738
transform 1 0 68 0 1 3
box -6 -4 34 96
use and2_1x  and2_1x_2
timestamp 1484419738
transform 1 0 100 0 1 3
box -6 -4 34 96
use and2_1x  and2_1x_3
timestamp 1484419738
transform 1 0 132 0 1 3
box -6 -4 34 96
use and2_1x  and2_1x_4
timestamp 1484419738
transform 1 0 164 0 1 3
box -6 -4 34 96
use and2_1x  and2_1x_5
timestamp 1484419738
transform 1 0 196 0 1 3
box -6 -4 34 96
use and2_1x  and2_1x_6
timestamp 1484419738
transform 1 0 228 0 1 3
box -6 -4 34 96
use inv_1x  inv_1x_0
timestamp 1484418501
transform 1 0 -316 0 1 -127
box -6 -4 18 96
use and2_1x  and2_1x_7
timestamp 1484419738
transform 1 0 -300 0 1 -127
box -6 -4 34 96
use mux2_dp_1x  mux2_dp_1x_20
timestamp 1484435125
transform 1 0 -268 0 1 -127
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_17
timestamp 1484435125
transform 1 0 -220 0 1 -127
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_16
timestamp 1484435125
transform 1 0 -172 0 1 -127
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_15
timestamp 1484435125
transform 1 0 -124 0 1 -127
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_14
timestamp 1484435125
transform 1 0 -76 0 1 -127
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_13
timestamp 1484435125
transform 1 0 -28 0 1 -127
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_12
timestamp 1484435125
transform 1 0 20 0 1 -127
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_11
timestamp 1484435125
transform 1 0 68 0 1 -127
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_10
timestamp 1484435125
transform 1 0 116 0 1 -127
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_9
timestamp 1484435125
transform 1 0 164 0 1 -127
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_8
timestamp 1484435125
transform 1 0 212 0 1 -127
box -6 -4 50 96
use xor2_1x  xor2_1x_0
timestamp 1492273518
transform 1 0 -228 0 1 -257
box -6 -4 58 96
use mux2_dp_1x  mux2_dp_1x_27
timestamp 1484435125
transform 1 0 -172 0 1 -257
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_26
timestamp 1484435125
transform 1 0 -124 0 1 -257
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_25
timestamp 1484435125
transform 1 0 -76 0 1 -257
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_24
timestamp 1484435125
transform 1 0 -28 0 1 -257
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_23
timestamp 1484435125
transform 1 0 20 0 1 -257
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_22
timestamp 1484435125
transform 1 0 68 0 1 -257
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_21
timestamp 1484435125
transform 1 0 116 0 1 -257
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_19
timestamp 1484435125
transform 1 0 164 0 1 -257
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_18
timestamp 1484435125
transform 1 0 212 0 1 -257
box -6 -4 50 96
use xor2_1x  xor2_1x_2
timestamp 1492273518
transform 1 0 -236 0 1 -387
box -6 -4 58 96
use xor2_1x  xor2_1x_1
timestamp 1492273518
transform 1 0 -180 0 1 -387
box -6 -4 58 96
use mux2_dp_1x  mux2_dp_1x_35
timestamp 1484435125
transform 1 0 -124 0 1 -387
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_34
timestamp 1484435125
transform 1 0 -76 0 1 -387
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_33
timestamp 1484435125
transform 1 0 -28 0 1 -387
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_32
timestamp 1484435125
transform 1 0 20 0 1 -387
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_31
timestamp 1484435125
transform 1 0 68 0 1 -387
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_30
timestamp 1484435125
transform 1 0 116 0 1 -387
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_29
timestamp 1484435125
transform 1 0 164 0 1 -387
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_28
timestamp 1484435125
transform 1 0 212 0 1 -387
box -6 -4 50 96
<< labels >>
rlabel metal1 -348 111 -348 111 1 a6
rlabel metal1 -348 118 -348 118 1 a5
rlabel metal1 -348 125 -348 125 1 a4
rlabel metal1 -348 132 -348 132 1 a3
rlabel metal1 -348 139 -348 139 1 a2
rlabel metal1 -348 146 -348 146 1 a1
rlabel metal1 -348 153 -348 153 5 a0
rlabel m3contact -328 -95 -328 -95 1 arith
rlabel metal3 -320 -18 -320 -18 1 right
rlabel metal3 -320 -27 -320 -27 1 rightb
rlabel metal3 -320 -9 -320 -9 1 arithAndRight
rlabel metal1 -348 104 -348 104 1 a7
<< end >>
